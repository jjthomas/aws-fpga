`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module DualPortBRAM(
  input         clock,
  input  [4:0]  io_a_addr,
  input  [15:0] io_a_din,
  input         io_a_wr,
  input  [4:0]  io_b_addr,
  output [15:0] io_b_dout
);
  reg [15:0] mem [0:31];
  reg [31:0] _RAND_0;
  wire [15:0] mem__T_12_data;
  wire [4:0] mem__T_12_addr;
  wire [15:0] mem__T_14_data;
  wire [4:0] mem__T_14_addr;
  wire [15:0] mem__T_13_data;
  wire [4:0] mem__T_13_addr;
  wire  mem__T_13_mask;
  wire  mem__T_13_en;
  wire [15:0] mem__T_15_data;
  wire [4:0] mem__T_15_addr;
  wire  mem__T_15_mask;
  wire  mem__T_15_en;
  wire  _GEN_8;
  reg [4:0] mem__T_12_addr_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] mem__T_14_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign mem__T_12_addr = mem__T_12_addr_pipe_0;
  assign mem__T_12_data = mem[mem__T_12_addr];
  assign mem__T_14_addr = mem__T_14_addr_pipe_0;
  assign mem__T_14_data = mem[mem__T_14_addr];
  assign mem__T_13_data = io_a_din;
  assign mem__T_13_addr = io_a_addr;
  assign mem__T_13_mask = io_a_wr;
  assign mem__T_13_en = io_a_wr;
  assign mem__T_15_data = 16'h0;
  assign mem__T_15_addr = io_b_addr;
  assign mem__T_15_mask = 1'h0;
  assign mem__T_15_en = 1'h0;
  assign _GEN_8 = 1'h1;
  assign io_b_dout = mem__T_14_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem__T_12_addr_pipe_0 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem__T_14_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_13_en & mem__T_13_mask) begin
      mem[mem__T_13_addr] <= mem__T_13_data;
    end
    if(mem__T_15_en & mem__T_15_mask) begin
      mem[mem__T_15_addr] <= mem__T_15_data;
    end
    if (_GEN_8) begin
      mem__T_12_addr_pipe_0 <= io_a_addr;
    end
    if (_GEN_8) begin
      mem__T_14_addr_pipe_0 <= io_b_addr;
    end
  end
endmodule
module PassThrough(
  input         clock,
  input         reset,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  input  [9:0]  io_inputBits,
  output        io_inputMemConsumed,
  input         io_inputFinished,
  output [15:0] io_outputMemBlock,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output [9:0]  io_outputBits,
  output        io_outputFinished,
  input         io_outputMemFlushed
);
  reg  inputMemBlock_0;
  reg [31:0] _RAND_0;
  reg  inputMemBlock_1;
  reg [31:0] _RAND_1;
  reg  inputMemBlock_2;
  reg [31:0] _RAND_2;
  reg  inputMemBlock_3;
  reg [31:0] _RAND_3;
  reg  inputMemBlock_4;
  reg [31:0] _RAND_4;
  reg  inputMemBlock_5;
  reg [31:0] _RAND_5;
  reg  inputMemBlock_6;
  reg [31:0] _RAND_6;
  reg  inputMemBlock_7;
  reg [31:0] _RAND_7;
  reg  inputMemBlock_8;
  reg [31:0] _RAND_8;
  reg  inputMemBlock_9;
  reg [31:0] _RAND_9;
  reg  inputMemBlock_10;
  reg [31:0] _RAND_10;
  reg  inputMemBlock_11;
  reg [31:0] _RAND_11;
  reg  inputMemBlock_12;
  reg [31:0] _RAND_12;
  reg  inputMemBlock_13;
  reg [31:0] _RAND_13;
  reg  inputMemBlock_14;
  reg [31:0] _RAND_14;
  reg  inputMemBlock_15;
  reg [31:0] _RAND_15;
  reg [4:0] inputPieceBitsRemaining;
  reg [31:0] _RAND_16;
  reg [9:0] inputBitsRemaining;
  reg [31:0] _RAND_17;
  reg  inputBlockLoaded;
  reg [31:0] _RAND_18;
  reg  outputMemBlock_0;
  reg [31:0] _RAND_19;
  reg  outputMemBlock_1;
  reg [31:0] _RAND_20;
  reg  outputMemBlock_2;
  reg [31:0] _RAND_21;
  reg  outputMemBlock_3;
  reg [31:0] _RAND_22;
  reg  outputMemBlock_4;
  reg [31:0] _RAND_23;
  reg  outputMemBlock_5;
  reg [31:0] _RAND_24;
  reg  outputMemBlock_6;
  reg [31:0] _RAND_25;
  reg  outputMemBlock_7;
  reg [31:0] _RAND_26;
  reg  outputMemBlock_8;
  reg [31:0] _RAND_27;
  reg  outputMemBlock_9;
  reg [31:0] _RAND_28;
  reg  outputMemBlock_10;
  reg [31:0] _RAND_29;
  reg  outputMemBlock_11;
  reg [31:0] _RAND_30;
  reg  outputMemBlock_12;
  reg [31:0] _RAND_31;
  reg  outputMemBlock_13;
  reg [31:0] _RAND_32;
  reg  outputMemBlock_14;
  reg [31:0] _RAND_33;
  reg  outputMemBlock_15;
  reg [31:0] _RAND_34;
  reg [9:0] outputBits;
  reg [31:0] _RAND_35;
  reg [4:0] outputPieceBits;
  reg [31:0] _RAND_36;
  wire  inputBram_clock;
  wire [4:0] inputBram_io_a_addr;
  wire [15:0] inputBram_io_a_din;
  wire  inputBram_io_a_wr;
  wire [4:0] inputBram_io_b_addr;
  wire [15:0] inputBram_io_b_dout;
  reg [4:0] inputReadAddr;
  reg [31:0] _RAND_37;
  reg  inputPieceRead;
  reg [31:0] _RAND_38;
  wire  outputBram_clock;
  wire [4:0] outputBram_io_a_addr;
  wire [15:0] outputBram_io_a_din;
  wire  outputBram_io_a_wr;
  wire [4:0] outputBram_io_b_addr;
  wire [15:0] outputBram_io_b_dout;
  reg [4:0] outputWriteAddr;
  reg [31:0] _RAND_39;
  reg [4:0] outputReadAddr;
  reg [31:0] _RAND_40;
  wire  _T_75;
  wire  _T_76;
  wire  _GEN_0;
  wire [9:0] _GEN_1;
  wire  _T_79;
  wire  _T_80;
  wire  _GEN_2;
  wire  _T_84;
  wire  _T_85;
  wire  _T_87;
  wire  _T_88;
  wire  _T_90;
  wire  _T_94;
  wire [9:0] _T_96;
  wire [5:0] _T_98;
  wire [4:0] _T_99;
  wire  _T_100;
  wire  _T_101;
  wire  _T_102;
  wire  _T_103;
  wire  _T_104;
  wire  _T_105;
  wire  _T_106;
  wire  _T_107;
  wire  _T_108;
  wire  _T_109;
  wire  _T_110;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  _T_114;
  wire  _T_115;
  wire [9:0] _GEN_4;
  wire [4:0] _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [9:0] _GEN_23;
  wire [4:0] _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  inputAdvance;
  wire  _T_118;
  wire  _T_120;
  wire  _T_122;
  wire  _T_123;
  wire  _T_125;
  wire  _T_126;
  wire [5:0] _T_128;
  wire [5:0] _T_129;
  wire [4:0] _T_130;
  wire [10:0] _T_132;
  wire [10:0] _T_133;
  wire [9:0] _T_134;
  wire [9:0] _GEN_41;
  wire [9:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  nextBitValid;
  wire  nextBit;
  wire [5:0] _T_138;
  wire [4:0] _T_139;
  wire [10:0] _T_141;
  wire [9:0] _T_142;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire [4:0] _GEN_74;
  wire [9:0] _GEN_75;
  wire  _T_144;
  wire  _T_147;
  wire  _T_149;
  wire  _T_150;
  wire  _T_151;
  wire [1:0] _T_152;
  wire [1:0] _T_153;
  wire [3:0] _T_154;
  wire [1:0] _T_155;
  wire [1:0] _T_156;
  wire [3:0] _T_157;
  wire [7:0] _T_158;
  wire [1:0] _T_159;
  wire [1:0] _T_160;
  wire [3:0] _T_161;
  wire [1:0] _T_162;
  wire [1:0] _T_163;
  wire [3:0] _T_164;
  wire [7:0] _T_165;
  wire [15:0] _T_166;
  wire [5:0] _T_171;
  wire [4:0] _T_172;
  wire [4:0] _GEN_76;
  wire [4:0] _GEN_77;
  reg  outputReadingStarted;
  reg [31:0] _RAND_41;
  wire  _T_177;
  wire  _T_184;
  wire  _T_185;
  wire  _T_186;
  wire  _T_187;
  wire  _GEN_78;
  wire  _T_189;
  wire  _T_191;
  wire  _T_192;
  wire [5:0] _T_194;
  wire [4:0] _T_195;
  wire [4:0] _GEN_79;
  wire  _T_199;
  wire  _T_200;
  wire  _T_210;
  wire  _T_215;
  wire  _T_216;
  wire [9:0] _GEN_80;
  wire [4:0] _GEN_81;
  wire  _GEN_82;
  wire [4:0] _GEN_83;
  wire [4:0] _GEN_84;
  DualPortBRAM inputBram (
    .clock(inputBram_clock),
    .io_a_addr(inputBram_io_a_addr),
    .io_a_din(inputBram_io_a_din),
    .io_a_wr(inputBram_io_a_wr),
    .io_b_addr(inputBram_io_b_addr),
    .io_b_dout(inputBram_io_b_dout)
  );
  DualPortBRAM outputBram (
    .clock(outputBram_clock),
    .io_a_addr(outputBram_io_a_addr),
    .io_a_din(outputBram_io_a_din),
    .io_a_wr(outputBram_io_a_wr),
    .io_b_addr(outputBram_io_b_addr),
    .io_b_dout(outputBram_io_b_dout)
  );
  assign _T_75 = io_inputMemIdx == 5'h1f;
  assign _T_76 = io_inputMemBlockValid & _T_75;
  assign _GEN_0 = _T_76 ? 1'h1 : inputBlockLoaded;
  assign _GEN_1 = _T_76 ? io_inputBits : inputBitsRemaining;
  assign _T_79 = inputBitsRemaining == 10'h0;
  assign _T_80 = inputBlockLoaded & _T_79;
  assign _GEN_2 = _T_80 ? 1'h0 : _GEN_0;
  assign _T_84 = inputPieceBitsRemaining == 5'h0;
  assign _T_85 = inputBlockLoaded & _T_84;
  assign _T_87 = inputBitsRemaining != 10'h0;
  assign _T_88 = _T_85 & _T_87;
  assign _T_90 = inputPieceRead == 1'h0;
  assign _T_94 = inputBitsRemaining < 10'h10;
  assign _T_96 = _T_94 ? inputBitsRemaining : 10'h10;
  assign _T_98 = inputReadAddr + 5'h1;
  assign _T_99 = _T_98[4:0];
  assign _T_100 = inputBram_io_b_dout[0];
  assign _T_101 = inputBram_io_b_dout[1];
  assign _T_102 = inputBram_io_b_dout[2];
  assign _T_103 = inputBram_io_b_dout[3];
  assign _T_104 = inputBram_io_b_dout[4];
  assign _T_105 = inputBram_io_b_dout[5];
  assign _T_106 = inputBram_io_b_dout[6];
  assign _T_107 = inputBram_io_b_dout[7];
  assign _T_108 = inputBram_io_b_dout[8];
  assign _T_109 = inputBram_io_b_dout[9];
  assign _T_110 = inputBram_io_b_dout[10];
  assign _T_111 = inputBram_io_b_dout[11];
  assign _T_112 = inputBram_io_b_dout[12];
  assign _T_113 = inputBram_io_b_dout[13];
  assign _T_114 = inputBram_io_b_dout[14];
  assign _T_115 = inputBram_io_b_dout[15];
  assign _GEN_4 = _T_90 ? {{5'd0}, inputPieceBitsRemaining} : _T_96;
  assign _GEN_5 = _T_90 ? inputReadAddr : _T_99;
  assign _GEN_6 = _T_90 ? inputMemBlock_0 : _T_100;
  assign _GEN_7 = _T_90 ? inputMemBlock_1 : _T_101;
  assign _GEN_8 = _T_90 ? inputMemBlock_2 : _T_102;
  assign _GEN_9 = _T_90 ? inputMemBlock_3 : _T_103;
  assign _GEN_10 = _T_90 ? inputMemBlock_4 : _T_104;
  assign _GEN_11 = _T_90 ? inputMemBlock_5 : _T_105;
  assign _GEN_12 = _T_90 ? inputMemBlock_6 : _T_106;
  assign _GEN_13 = _T_90 ? inputMemBlock_7 : _T_107;
  assign _GEN_14 = _T_90 ? inputMemBlock_8 : _T_108;
  assign _GEN_15 = _T_90 ? inputMemBlock_9 : _T_109;
  assign _GEN_16 = _T_90 ? inputMemBlock_10 : _T_110;
  assign _GEN_17 = _T_90 ? inputMemBlock_11 : _T_111;
  assign _GEN_18 = _T_90 ? inputMemBlock_12 : _T_112;
  assign _GEN_19 = _T_90 ? inputMemBlock_13 : _T_113;
  assign _GEN_20 = _T_90 ? inputMemBlock_14 : _T_114;
  assign _GEN_21 = _T_90 ? inputMemBlock_15 : _T_115;
  assign _GEN_22 = _T_88 ? _T_90 : inputPieceRead;
  assign _GEN_23 = _T_88 ? _GEN_4 : {{5'd0}, inputPieceBitsRemaining};
  assign _GEN_24 = _T_88 ? _GEN_5 : inputReadAddr;
  assign _GEN_25 = _T_88 ? _GEN_6 : inputMemBlock_0;
  assign _GEN_26 = _T_88 ? _GEN_7 : inputMemBlock_1;
  assign _GEN_27 = _T_88 ? _GEN_8 : inputMemBlock_2;
  assign _GEN_28 = _T_88 ? _GEN_9 : inputMemBlock_3;
  assign _GEN_29 = _T_88 ? _GEN_10 : inputMemBlock_4;
  assign _GEN_30 = _T_88 ? _GEN_11 : inputMemBlock_5;
  assign _GEN_31 = _T_88 ? _GEN_12 : inputMemBlock_6;
  assign _GEN_32 = _T_88 ? _GEN_13 : inputMemBlock_7;
  assign _GEN_33 = _T_88 ? _GEN_14 : inputMemBlock_8;
  assign _GEN_34 = _T_88 ? _GEN_15 : inputMemBlock_9;
  assign _GEN_35 = _T_88 ? _GEN_16 : inputMemBlock_10;
  assign _GEN_36 = _T_88 ? _GEN_17 : inputMemBlock_11;
  assign _GEN_37 = _T_88 ? _GEN_18 : inputMemBlock_12;
  assign _GEN_38 = _T_88 ? _GEN_19 : inputMemBlock_13;
  assign _GEN_39 = _T_88 ? _GEN_20 : inputMemBlock_14;
  assign _GEN_40 = _T_88 ? _GEN_21 : inputMemBlock_15;
  assign _T_118 = outputPieceBits != 5'h10;
  assign _T_120 = outputBits == 10'h200;
  assign _T_122 = _T_120 == 1'h0;
  assign _T_123 = _T_118 & _T_122;
  assign _T_125 = inputPieceBitsRemaining != 5'h0;
  assign _T_126 = _T_123 & _T_125;
  assign _T_128 = inputPieceBitsRemaining - 5'h1;
  assign _T_129 = $unsigned(_T_128);
  assign _T_130 = _T_129[4:0];
  assign _T_132 = inputBitsRemaining - 10'h1;
  assign _T_133 = $unsigned(_T_132);
  assign _T_134 = _T_133[9:0];
  assign _GEN_41 = inputAdvance ? {{5'd0}, _T_130} : _GEN_23;
  assign _GEN_42 = inputAdvance ? _T_134 : _GEN_1;
  assign _GEN_43 = inputAdvance ? inputMemBlock_1 : _GEN_25;
  assign _GEN_44 = inputAdvance ? inputMemBlock_2 : _GEN_26;
  assign _GEN_45 = inputAdvance ? inputMemBlock_3 : _GEN_27;
  assign _GEN_46 = inputAdvance ? inputMemBlock_4 : _GEN_28;
  assign _GEN_47 = inputAdvance ? inputMemBlock_5 : _GEN_29;
  assign _GEN_48 = inputAdvance ? inputMemBlock_6 : _GEN_30;
  assign _GEN_49 = inputAdvance ? inputMemBlock_7 : _GEN_31;
  assign _GEN_50 = inputAdvance ? inputMemBlock_8 : _GEN_32;
  assign _GEN_51 = inputAdvance ? inputMemBlock_9 : _GEN_33;
  assign _GEN_52 = inputAdvance ? inputMemBlock_10 : _GEN_34;
  assign _GEN_53 = inputAdvance ? inputMemBlock_11 : _GEN_35;
  assign _GEN_54 = inputAdvance ? inputMemBlock_12 : _GEN_36;
  assign _GEN_55 = inputAdvance ? inputMemBlock_13 : _GEN_37;
  assign _GEN_56 = inputAdvance ? inputMemBlock_14 : _GEN_38;
  assign _GEN_57 = inputAdvance ? inputMemBlock_15 : _GEN_39;
  assign _T_138 = outputPieceBits + 5'h1;
  assign _T_139 = _T_138[4:0];
  assign _T_141 = outputBits + 10'h1;
  assign _T_142 = _T_141[9:0];
  assign _GEN_58 = nextBitValid ? nextBit : outputMemBlock_15;
  assign _GEN_59 = nextBitValid ? outputMemBlock_1 : outputMemBlock_0;
  assign _GEN_60 = nextBitValid ? outputMemBlock_2 : outputMemBlock_1;
  assign _GEN_61 = nextBitValid ? outputMemBlock_3 : outputMemBlock_2;
  assign _GEN_62 = nextBitValid ? outputMemBlock_4 : outputMemBlock_3;
  assign _GEN_63 = nextBitValid ? outputMemBlock_5 : outputMemBlock_4;
  assign _GEN_64 = nextBitValid ? outputMemBlock_6 : outputMemBlock_5;
  assign _GEN_65 = nextBitValid ? outputMemBlock_7 : outputMemBlock_6;
  assign _GEN_66 = nextBitValid ? outputMemBlock_8 : outputMemBlock_7;
  assign _GEN_67 = nextBitValid ? outputMemBlock_9 : outputMemBlock_8;
  assign _GEN_68 = nextBitValid ? outputMemBlock_10 : outputMemBlock_9;
  assign _GEN_69 = nextBitValid ? outputMemBlock_11 : outputMemBlock_10;
  assign _GEN_70 = nextBitValid ? outputMemBlock_12 : outputMemBlock_11;
  assign _GEN_71 = nextBitValid ? outputMemBlock_13 : outputMemBlock_12;
  assign _GEN_72 = nextBitValid ? outputMemBlock_14 : outputMemBlock_13;
  assign _GEN_73 = nextBitValid ? outputMemBlock_15 : outputMemBlock_14;
  assign _GEN_74 = nextBitValid ? _T_139 : outputPieceBits;
  assign _GEN_75 = nextBitValid ? _T_142 : outputBits;
  assign _T_144 = outputPieceBits == 5'h10;
  assign _T_147 = io_inputFinished & _T_79;
  assign _T_149 = outputPieceBits > 5'h0;
  assign _T_150 = _T_147 & _T_149;
  assign _T_151 = _T_144 | _T_150;
  assign _T_152 = {outputMemBlock_1,outputMemBlock_0};
  assign _T_153 = {outputMemBlock_3,outputMemBlock_2};
  assign _T_154 = {_T_153,_T_152};
  assign _T_155 = {outputMemBlock_5,outputMemBlock_4};
  assign _T_156 = {outputMemBlock_7,outputMemBlock_6};
  assign _T_157 = {_T_156,_T_155};
  assign _T_158 = {_T_157,_T_154};
  assign _T_159 = {outputMemBlock_9,outputMemBlock_8};
  assign _T_160 = {outputMemBlock_11,outputMemBlock_10};
  assign _T_161 = {_T_160,_T_159};
  assign _T_162 = {outputMemBlock_13,outputMemBlock_12};
  assign _T_163 = {outputMemBlock_15,outputMemBlock_14};
  assign _T_164 = {_T_163,_T_162};
  assign _T_165 = {_T_164,_T_161};
  assign _T_166 = {_T_165,_T_158};
  assign _T_171 = outputWriteAddr + 5'h1;
  assign _T_172 = _T_171[4:0];
  assign _GEN_76 = _T_144 ? 5'h0 : _GEN_74;
  assign _GEN_77 = _T_144 ? _T_172 : outputWriteAddr;
  assign _T_177 = outputReadingStarted == 1'h0;
  assign _T_184 = outputBits > 10'h0;
  assign _T_185 = _T_147 & _T_184;
  assign _T_186 = _T_120 | _T_185;
  assign _T_187 = _T_177 & _T_186;
  assign _GEN_78 = _T_187 ? 1'h1 : outputReadingStarted;
  assign _T_189 = io_outputMemBlockReady & outputReadingStarted;
  assign _T_191 = outputReadAddr != 5'h1f;
  assign _T_192 = _T_189 & _T_191;
  assign _T_194 = outputReadAddr + 5'h1;
  assign _T_195 = _T_194[4:0];
  assign _GEN_79 = _T_192 ? _T_195 : outputReadAddr;
  assign _T_199 = io_inputFinished == 1'h0;
  assign _T_200 = _T_79 & _T_199;
  assign _T_210 = outputReadingStarted & _T_186;
  assign _T_215 = outputBits == 10'h0;
  assign _T_216 = _T_147 & _T_215;
  assign _GEN_80 = io_outputMemFlushed ? 10'h0 : _GEN_75;
  assign _GEN_81 = io_outputMemFlushed ? 5'h0 : _GEN_76;
  assign _GEN_82 = io_outputMemFlushed ? 1'h0 : _GEN_78;
  assign _GEN_83 = io_outputMemFlushed ? 5'h0 : _GEN_77;
  assign _GEN_84 = io_outputMemFlushed ? 5'h0 : _GEN_79;
  assign io_inputMemConsumed = _T_200;
  assign io_outputMemBlock = outputBram_io_b_dout;
  assign io_outputMemBlockValid = _T_210;
  assign io_outputBits = outputBits;
  assign io_outputFinished = _T_216;
  assign inputBram_io_a_addr = io_inputMemIdx;
  assign inputBram_io_a_din = io_inputMemBlock;
  assign inputBram_io_a_wr = io_inputMemBlockValid;
  assign inputBram_io_b_addr = inputReadAddr;
  assign inputBram_clock = clock;
  assign outputBram_io_a_addr = outputWriteAddr;
  assign outputBram_io_a_din = _T_166;
  assign outputBram_io_a_wr = _T_151;
  assign outputBram_io_b_addr = outputReadAddr;
  assign outputBram_clock = clock;
  assign inputAdvance = _T_126;
  assign nextBitValid = inputAdvance;
  assign nextBit = inputMemBlock_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  inputMemBlock_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  inputMemBlock_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputMemBlock_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  inputMemBlock_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  inputMemBlock_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  inputMemBlock_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  inputMemBlock_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemBlock_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBlock_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  inputMemBlock_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputMemBlock_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  inputMemBlock_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  inputMemBlock_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  inputMemBlock_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  inputMemBlock_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  inputMemBlock_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  inputPieceBitsRemaining = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  inputBitsRemaining = _RAND_17[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  inputBlockLoaded = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  outputMemBlock_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  outputMemBlock_1 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  outputMemBlock_2 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  outputMemBlock_3 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  outputMemBlock_4 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  outputMemBlock_5 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  outputMemBlock_6 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  outputMemBlock_7 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  outputMemBlock_8 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  outputMemBlock_9 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  outputMemBlock_10 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  outputMemBlock_11 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  outputMemBlock_12 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  outputMemBlock_13 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  outputMemBlock_14 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  outputMemBlock_15 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  outputBits = _RAND_35[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  outputPieceBits = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  inputReadAddr = _RAND_37[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  inputPieceRead = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  outputWriteAddr = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  outputReadAddr = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  outputReadingStarted = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (inputAdvance) begin
      inputMemBlock_0 <= inputMemBlock_1;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_0 <= _T_100;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_1 <= inputMemBlock_2;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_1 <= _T_101;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_2 <= inputMemBlock_3;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_2 <= _T_102;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_3 <= inputMemBlock_4;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_3 <= _T_103;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_4 <= inputMemBlock_5;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_4 <= _T_104;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_5 <= inputMemBlock_6;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_5 <= _T_105;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_6 <= inputMemBlock_7;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_6 <= _T_106;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_7 <= inputMemBlock_8;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_7 <= _T_107;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_8 <= inputMemBlock_9;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_8 <= _T_108;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_9 <= inputMemBlock_10;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_9 <= _T_109;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_10 <= inputMemBlock_11;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_10 <= _T_110;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_11 <= inputMemBlock_12;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_11 <= _T_111;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_12 <= inputMemBlock_13;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_12 <= _T_112;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_13 <= inputMemBlock_14;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_13 <= _T_113;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_14 <= inputMemBlock_15;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_14 <= _T_114;
        end
      end
    end
    if (_T_88) begin
      if (!(_T_90)) begin
        inputMemBlock_15 <= _T_115;
      end
    end
    if (reset) begin
      inputPieceBitsRemaining <= 5'h0;
    end else begin
      inputPieceBitsRemaining <= _GEN_41[4:0];
    end
    if (reset) begin
      inputBitsRemaining <= 10'h0;
    end else begin
      if (inputAdvance) begin
        inputBitsRemaining <= _T_134;
      end else begin
        if (_T_76) begin
          inputBitsRemaining <= io_inputBits;
        end
      end
    end
    if (reset) begin
      inputBlockLoaded <= 1'h0;
    end else begin
      if (_T_80) begin
        inputBlockLoaded <= 1'h0;
      end else begin
        if (_T_76) begin
          inputBlockLoaded <= 1'h1;
        end
      end
    end
    if (nextBitValid) begin
      outputMemBlock_0 <= outputMemBlock_1;
    end
    if (nextBitValid) begin
      outputMemBlock_1 <= outputMemBlock_2;
    end
    if (nextBitValid) begin
      outputMemBlock_2 <= outputMemBlock_3;
    end
    if (nextBitValid) begin
      outputMemBlock_3 <= outputMemBlock_4;
    end
    if (nextBitValid) begin
      outputMemBlock_4 <= outputMemBlock_5;
    end
    if (nextBitValid) begin
      outputMemBlock_5 <= outputMemBlock_6;
    end
    if (nextBitValid) begin
      outputMemBlock_6 <= outputMemBlock_7;
    end
    if (nextBitValid) begin
      outputMemBlock_7 <= outputMemBlock_8;
    end
    if (nextBitValid) begin
      outputMemBlock_8 <= outputMemBlock_9;
    end
    if (nextBitValid) begin
      outputMemBlock_9 <= outputMemBlock_10;
    end
    if (nextBitValid) begin
      outputMemBlock_10 <= outputMemBlock_11;
    end
    if (nextBitValid) begin
      outputMemBlock_11 <= outputMemBlock_12;
    end
    if (nextBitValid) begin
      outputMemBlock_12 <= outputMemBlock_13;
    end
    if (nextBitValid) begin
      outputMemBlock_13 <= outputMemBlock_14;
    end
    if (nextBitValid) begin
      outputMemBlock_14 <= outputMemBlock_15;
    end
    if (nextBitValid) begin
      outputMemBlock_15 <= nextBit;
    end
    if (reset) begin
      outputBits <= 10'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputBits <= 10'h0;
      end else begin
        if (nextBitValid) begin
          outputBits <= _T_142;
        end
      end
    end
    if (reset) begin
      outputPieceBits <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputPieceBits <= 5'h0;
      end else begin
        if (_T_144) begin
          outputPieceBits <= 5'h0;
        end else begin
          if (nextBitValid) begin
            outputPieceBits <= _T_139;
          end
        end
      end
    end
    if (reset) begin
      inputReadAddr <= 5'h0;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputReadAddr <= _T_99;
        end
      end
    end
    if (reset) begin
      inputPieceRead <= 1'h0;
    end else begin
      if (_T_88) begin
        inputPieceRead <= _T_90;
      end
    end
    if (reset) begin
      outputWriteAddr <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputWriteAddr <= 5'h0;
      end else begin
        if (_T_144) begin
          outputWriteAddr <= _T_172;
        end
      end
    end
    if (reset) begin
      outputReadAddr <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputReadAddr <= 5'h0;
      end else begin
        if (_T_192) begin
          outputReadAddr <= _T_195;
        end
      end
    end
    if (reset) begin
      outputReadingStarted <= 1'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputReadingStarted <= 1'h0;
      end else begin
        if (_T_187) begin
          outputReadingStarted <= 1'h1;
        end
      end
    end
  end
endmodule
module StreamingCore(
  input         clock,
  input         reset,
  output [63:0] io_inputMemAddr,
  output        io_inputMemAddrValid,
  input         io_inputMemAddrReady,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output        io_inputMemBlockReady,
  output [63:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [15:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output        io_inputFinished,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [15:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [15:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [63:0] inputBitsRemaining;
  reg [63:0] _RAND_2;
  reg  coreInputFinished;
  reg [31:0] _RAND_3;
  reg [63:0] outputBits;
  reg [63:0] _RAND_4;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_5;
  reg  outputLengthCommitted;
  reg [31:0] _RAND_6;
  reg [63:0] inputMemAddr;
  reg [63:0] _RAND_7;
  reg [63:0] outputMemAddr;
  reg [63:0] _RAND_8;
  reg [63:0] outputLenAddr;
  reg [63:0] _RAND_9;
  reg  inputAddressAccepted;
  reg [31:0] _RAND_10;
  wire  _T_41;
  wire  _T_42;
  wire  _T_44;
  wire  _T_46;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_53;
  wire  _GEN_0;
  wire  inputBlockReadable;
  wire  _T_56;
  wire  _T_57;
  wire  _T_59;
  wire [9:0] _T_61;
  wire [9:0] _T_62;
  wire  _T_64;
  wire [47:0] _T_65;
  wire [63:0] _T_66;
  wire [63:0] _GEN_1;
  wire  _T_68;
  wire [31:0] _T_69;
  wire [47:0] _T_70;
  wire [15:0] _T_71;
  wire [63:0] _T_72;
  wire [63:0] _GEN_2;
  wire  _T_74;
  wire [15:0] _T_75;
  wire [31:0] _T_76;
  wire [31:0] _T_77;
  wire [63:0] _T_78;
  wire [63:0] _GEN_3;
  wire  _T_80;
  wire [47:0] _T_81;
  wire [63:0] _T_82;
  wire [63:0] _GEN_4;
  wire  _T_84;
  wire [47:0] _T_85;
  wire [63:0] _T_86;
  wire [63:0] _GEN_5;
  wire  _T_88;
  wire [31:0] _T_89;
  wire [47:0] _T_90;
  wire [15:0] _T_91;
  wire [63:0] _T_92;
  wire [63:0] _GEN_6;
  wire  _T_94;
  wire [15:0] _T_95;
  wire [31:0] _T_96;
  wire [31:0] _T_97;
  wire [63:0] _T_98;
  wire [63:0] _GEN_7;
  wire  _T_100;
  wire [47:0] _T_101;
  wire [63:0] _T_102;
  wire [63:0] _GEN_8;
  wire  _T_104;
  wire [47:0] _T_105;
  wire [63:0] _T_106;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire  _T_108;
  wire [31:0] _T_109;
  wire [47:0] _T_110;
  wire [15:0] _T_111;
  wire [63:0] _T_112;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire  _T_114;
  wire [15:0] _T_115;
  wire [31:0] _T_116;
  wire [31:0] _T_117;
  wire [63:0] _T_118;
  wire [63:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire  _T_120;
  wire [47:0] _T_121;
  wire [63:0] _T_122;
  wire [63:0] _GEN_15;
  wire [63:0] _GEN_16;
  wire  _T_124;
  wire [64:0] _T_128;
  wire [63:0] _T_129;
  wire  _GEN_17;
  wire  _GEN_18;
  wire [63:0] _GEN_19;
  wire [64:0] _T_135;
  wire [64:0] _T_136;
  wire [63:0] _T_137;
  wire [63:0] _T_139;
  wire [64:0] _T_141;
  wire [63:0] _T_142;
  wire [63:0] _GEN_20;
  wire [63:0] _GEN_21;
  wire [63:0] _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [63:0] _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire [63:0] _GEN_29;
  wire [63:0] _GEN_30;
  wire [63:0] _GEN_31;
  wire [63:0] _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _T_150;
  wire  _GEN_36;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_11;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_12;
  wire  _GEN_37;
  wire [63:0] _T_157;
  wire  _T_159;
  wire  _T_161;
  wire  _T_162;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _GEN_38;
  wire  _T_171;
  wire [4:0] _GEN_39;
  wire [5:0] _T_174;
  wire [4:0] _T_175;
  wire [4:0] _GEN_40;
  wire [4:0] _GEN_41;
  wire [15:0] outputBitsBlock;
  wire  _T_178;
  wire [15:0] _T_179;
  wire  _T_181;
  wire [15:0] _T_182;
  wire  _T_184;
  wire [15:0] _T_185;
  wire  _T_187;
  wire [15:0] _T_188;
  wire [15:0] _T_190;
  wire [15:0] _T_191;
  wire [15:0] _T_192;
  wire [15:0] _T_193;
  wire [15:0] _T_194;
  wire  _T_195;
  wire  _T_199;
  wire [63:0] _GEN_50;
  wire [64:0] _T_203;
  wire [63:0] _T_204;
  wire  _GEN_42;
  wire [63:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire [63:0] _GEN_48;
  wire [63:0] _GEN_49;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign _T_41 = inputAddressAccepted == 1'h0;
  assign _T_42 = initDone & core_io_inputMemConsumed;
  assign _T_44 = inputBitsRemaining == 64'h0;
  assign _T_46 = _T_44 == 1'h0;
  assign _T_47 = _T_42 & _T_46;
  assign _T_48 = isInit | _T_47;
  assign _T_49 = _T_41 & _T_48;
  assign _T_50 = io_inputMemAddrValid & io_inputMemAddrReady;
  assign _T_53 = reset == 1'h0;
  assign _GEN_0 = _T_50 ? 1'h1 : inputAddressAccepted;
  assign _T_56 = inputAddressAccepted & io_inputMemBlockValid;
  assign _T_57 = inputBlockReadable & initDone;
  assign _T_59 = inputBitsRemaining > 64'h200;
  assign _T_61 = inputBitsRemaining[9:0];
  assign _T_62 = _T_59 ? 10'h200 : _T_61;
  assign _T_64 = io_inputMemIdx == 5'h0;
  assign _T_65 = inputMemAddr[63:16];
  assign _T_66 = {_T_65,io_inputMemBlock};
  assign _GEN_1 = _T_64 ? _T_66 : inputMemAddr;
  assign _T_68 = io_inputMemIdx == 5'h1;
  assign _T_69 = inputMemAddr[63:32];
  assign _T_70 = {_T_69,io_inputMemBlock};
  assign _T_71 = inputMemAddr[15:0];
  assign _T_72 = {_T_70,_T_71};
  assign _GEN_2 = _T_68 ? _T_72 : _GEN_1;
  assign _T_74 = io_inputMemIdx == 5'h2;
  assign _T_75 = inputMemAddr[63:48];
  assign _T_76 = {_T_75,io_inputMemBlock};
  assign _T_77 = inputMemAddr[31:0];
  assign _T_78 = {_T_76,_T_77};
  assign _GEN_3 = _T_74 ? _T_78 : _GEN_2;
  assign _T_80 = io_inputMemIdx == 5'h3;
  assign _T_81 = inputMemAddr[47:0];
  assign _T_82 = {io_inputMemBlock,_T_81};
  assign _GEN_4 = _T_80 ? _T_82 : _GEN_3;
  assign _T_84 = io_inputMemIdx == 5'h4;
  assign _T_85 = inputBitsRemaining[63:16];
  assign _T_86 = {_T_85,io_inputMemBlock};
  assign _GEN_5 = _T_84 ? _T_86 : inputBitsRemaining;
  assign _T_88 = io_inputMemIdx == 5'h5;
  assign _T_89 = inputBitsRemaining[63:32];
  assign _T_90 = {_T_89,io_inputMemBlock};
  assign _T_91 = inputBitsRemaining[15:0];
  assign _T_92 = {_T_90,_T_91};
  assign _GEN_6 = _T_88 ? _T_92 : _GEN_5;
  assign _T_94 = io_inputMemIdx == 5'h6;
  assign _T_95 = inputBitsRemaining[63:48];
  assign _T_96 = {_T_95,io_inputMemBlock};
  assign _T_97 = inputBitsRemaining[31:0];
  assign _T_98 = {_T_96,_T_97};
  assign _GEN_7 = _T_94 ? _T_98 : _GEN_6;
  assign _T_100 = io_inputMemIdx == 5'h7;
  assign _T_101 = inputBitsRemaining[47:0];
  assign _T_102 = {io_inputMemBlock,_T_101};
  assign _GEN_8 = _T_100 ? _T_102 : _GEN_7;
  assign _T_104 = io_inputMemIdx == 5'h8;
  assign _T_105 = outputMemAddr[63:16];
  assign _T_106 = {_T_105,io_inputMemBlock};
  assign _GEN_9 = _T_104 ? _T_106 : outputMemAddr;
  assign _GEN_10 = _T_104 ? _T_106 : outputLenAddr;
  assign _T_108 = io_inputMemIdx == 5'h9;
  assign _T_109 = outputMemAddr[63:32];
  assign _T_110 = {_T_109,io_inputMemBlock};
  assign _T_111 = outputMemAddr[15:0];
  assign _T_112 = {_T_110,_T_111};
  assign _GEN_11 = _T_108 ? _T_112 : _GEN_9;
  assign _GEN_12 = _T_108 ? _T_112 : _GEN_10;
  assign _T_114 = io_inputMemIdx == 5'ha;
  assign _T_115 = outputMemAddr[63:48];
  assign _T_116 = {_T_115,io_inputMemBlock};
  assign _T_117 = outputMemAddr[31:0];
  assign _T_118 = {_T_116,_T_117};
  assign _GEN_13 = _T_114 ? _T_118 : _GEN_11;
  assign _GEN_14 = _T_114 ? _T_118 : _GEN_12;
  assign _T_120 = io_inputMemIdx == 5'hb;
  assign _T_121 = outputMemAddr[47:0];
  assign _T_122 = {io_inputMemBlock,_T_121};
  assign _GEN_15 = _T_120 ? _T_122 : _GEN_13;
  assign _GEN_16 = _T_120 ? _T_122 : _GEN_14;
  assign _T_124 = io_inputMemIdx == 5'h1f;
  assign _T_128 = outputMemAddr + 64'h40;
  assign _T_129 = _T_128[63:0];
  assign _GEN_17 = _T_124 ? 1'h0 : isInit;
  assign _GEN_18 = _T_124 ? 1'h1 : initDone;
  assign _GEN_19 = _T_124 ? _T_129 : _GEN_15;
  assign _T_135 = inputBitsRemaining - 64'h200;
  assign _T_136 = $unsigned(_T_135);
  assign _T_137 = _T_136[63:0];
  assign _T_139 = _T_59 ? _T_137 : 64'h0;
  assign _T_141 = inputMemAddr + 64'h40;
  assign _T_142 = _T_141[63:0];
  assign _GEN_20 = _T_124 ? _T_139 : inputBitsRemaining;
  assign _GEN_21 = _T_124 ? _T_142 : inputMemAddr;
  assign _GEN_22 = isInit ? _GEN_4 : _GEN_21;
  assign _GEN_23 = isInit ? _GEN_8 : _GEN_20;
  assign _GEN_24 = isInit ? _GEN_19 : outputMemAddr;
  assign _GEN_25 = isInit ? _GEN_16 : outputLenAddr;
  assign _GEN_26 = isInit ? _GEN_17 : isInit;
  assign _GEN_27 = isInit ? _GEN_18 : initDone;
  assign _GEN_28 = _T_124 ? 1'h0 : _GEN_0;
  assign _GEN_29 = inputBlockReadable ? _GEN_22 : inputMemAddr;
  assign _GEN_30 = inputBlockReadable ? _GEN_23 : inputBitsRemaining;
  assign _GEN_31 = inputBlockReadable ? _GEN_24 : outputMemAddr;
  assign _GEN_32 = inputBlockReadable ? _GEN_25 : outputLenAddr;
  assign _GEN_33 = inputBlockReadable ? _GEN_26 : isInit;
  assign _GEN_34 = inputBlockReadable ? _GEN_27 : initDone;
  assign _GEN_35 = inputBlockReadable ? _GEN_28 : _GEN_0;
  assign _T_150 = core_io_inputMemConsumed & _T_44;
  assign _GEN_36 = _T_150 ? 1'h1 : coreInputFinished;
  assign _GEN_37 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_157 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_159 = outputAddressAccepted == 1'h0;
  assign _T_161 = outputLengthCommitted == 1'h0;
  assign _T_162 = core_io_outputFinished & _T_161;
  assign _T_163 = core_io_outputMemBlockValid | _T_162;
  assign _T_164 = _T_159 & _T_163;
  assign _T_165 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_38 = _T_165 ? 1'h1 : outputAddressAccepted;
  assign _T_171 = outputBlockCounter == 5'h1f;
  assign _GEN_39 = io_outputMemBlockReady ? 5'h0 : outputBlockCounter;
  assign _T_174 = outputBlockCounter + 5'h1;
  assign _T_175 = _T_174[4:0];
  assign _GEN_40 = _T_171 ? _GEN_39 : _T_175;
  assign _GEN_41 = outputAddressAcceptedNext ? _GEN_40 : outputBlockCounter;
  assign _T_178 = outputBlockCounter == 5'h0;
  assign _T_179 = outputBits[15:0];
  assign _T_181 = outputBlockCounter == 5'h1;
  assign _T_182 = outputBits[31:16];
  assign _T_184 = outputBlockCounter == 5'h2;
  assign _T_185 = outputBits[47:32];
  assign _T_187 = outputBlockCounter == 5'h3;
  assign _T_188 = outputBits[63:48];
  assign _T_190 = _T_187 ? _T_188 : 16'h0;
  assign _T_191 = _T_184 ? _T_185 : _T_190;
  assign _T_192 = _T_181 ? _T_182 : _T_191;
  assign _T_193 = _T_178 ? _T_179 : _T_192;
  assign _T_194 = core_io_outputFinished ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_195 = outputAddressAcceptedNext & io_outputMemBlockReady;
  assign _T_199 = _T_195 & _T_171;
  assign _GEN_50 = {{54'd0}, core_io_outputBits};
  assign _T_203 = outputBits + _GEN_50;
  assign _T_204 = _T_203[63:0];
  assign _GEN_42 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _GEN_43 = core_io_outputFinished ? outputBits : _T_204;
  assign _GEN_44 = core_io_outputFinished ? _GEN_31 : _T_129;
  assign _GEN_45 = _T_199 ? 1'h0 : _GEN_38;
  assign _GEN_46 = _T_199 ? 1'h0 : _GEN_37;
  assign _GEN_47 = _T_199 ? _GEN_42 : outputLengthCommitted;
  assign _GEN_48 = _T_199 ? _GEN_43 : outputBits;
  assign _GEN_49 = _T_199 ? _GEN_44 : _GEN_31;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemAddrValid = _T_49;
  assign io_inputMemBlockReady = inputAddressAccepted;
  assign io_outputMemAddr = _T_157;
  assign io_outputMemAddrValid = _T_164;
  assign io_outputMemBlock = _T_194;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_inputFinished = _T_44;
  assign io_outputFinished = outputLengthCommitted;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_57;
  assign core_io_inputBits = _T_62;
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_io_outputMemFlushed = _T_195;
  assign core_clock = clock;
  assign core_reset = reset;
  assign inputBlockReadable = _T_56;
  assign outputBitsBlock = _T_193;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{$random}};
  inputBitsRemaining = _RAND_2[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  coreInputFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{$random}};
  outputBits = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputBlockCounter = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputLengthCommitted = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{$random}};
  inputMemAddr = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{$random}};
  outputMemAddr = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{$random}};
  outputLenAddr = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputAddressAccepted = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  outputAddressAccepted = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  outputAddressAcceptedNext = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 64'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_100) begin
            inputBitsRemaining <= _T_102;
          end else begin
            if (_T_94) begin
              inputBitsRemaining <= _T_98;
            end else begin
              if (_T_88) begin
                inputBitsRemaining <= _T_92;
              end else begin
                if (_T_84) begin
                  inputBitsRemaining <= _T_86;
                end
              end
            end
          end
        end else begin
          if (_T_124) begin
            if (_T_59) begin
              inputBitsRemaining <= _T_137;
            end else begin
              inputBitsRemaining <= 64'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_150) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 64'h0;
    end else begin
      if (_T_199) begin
        if (!(core_io_outputFinished)) begin
          outputBits <= _T_204;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_171) begin
          if (io_outputMemBlockReady) begin
            outputBlockCounter <= 5'h0;
          end
        end else begin
          outputBlockCounter <= _T_175;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_199) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 64'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_80) begin
            inputMemAddr <= _T_82;
          end else begin
            if (_T_74) begin
              inputMemAddr <= _T_78;
            end else begin
              if (_T_68) begin
                inputMemAddr <= _T_72;
              end else begin
                if (_T_64) begin
                  inputMemAddr <= _T_66;
                end
              end
            end
          end
        end else begin
          if (_T_124) begin
            inputMemAddr <= _T_142;
          end
        end
      end
    end
    if (_T_199) begin
      if (core_io_outputFinished) begin
        if (inputBlockReadable) begin
          if (isInit) begin
            if (_T_124) begin
              outputMemAddr <= _T_129;
            end else begin
              if (_T_120) begin
                outputMemAddr <= _T_122;
              end else begin
                if (_T_114) begin
                  outputMemAddr <= _T_118;
                end else begin
                  if (_T_108) begin
                    outputMemAddr <= _T_112;
                  end else begin
                    if (_T_104) begin
                      outputMemAddr <= _T_106;
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        outputMemAddr <= _T_129;
      end
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            outputMemAddr <= _T_129;
          end else begin
            if (_T_120) begin
              outputMemAddr <= _T_122;
            end else begin
              if (_T_114) begin
                outputMemAddr <= _T_118;
              end else begin
                if (_T_108) begin
                  outputMemAddr <= _T_112;
                end else begin
                  if (_T_104) begin
                    outputMemAddr <= _T_106;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (inputBlockReadable) begin
      if (isInit) begin
        if (_T_120) begin
          outputLenAddr <= _T_122;
        end else begin
          if (_T_114) begin
            outputLenAddr <= _T_118;
          end else begin
            if (_T_108) begin
              outputLenAddr <= _T_112;
            end else begin
              if (_T_104) begin
                outputLenAddr <= _T_106;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      inputAddressAccepted <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (_T_124) begin
          inputAddressAccepted <= 1'h0;
        end else begin
          if (_T_50) begin
            inputAddressAccepted <= 1'h1;
          end
        end
      end else begin
        if (_T_50) begin
          inputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_199) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_165) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_199) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_50 & _T_53) begin
          $fwrite(32'h80000002,"input address 0x%h accepted for core 0\n",io_inputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_165 & _T_53) begin
          $fwrite(32'h80000002,"output address 0x%h accepted for core 0\n",io_outputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module StreamingCore_1(
  input         clock,
  input         reset,
  output [63:0] io_inputMemAddr,
  output        io_inputMemAddrValid,
  input         io_inputMemAddrReady,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output        io_inputMemBlockReady,
  output [63:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [15:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output        io_inputFinished,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [15:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [15:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [63:0] inputBitsRemaining;
  reg [63:0] _RAND_2;
  reg  coreInputFinished;
  reg [31:0] _RAND_3;
  reg [63:0] outputBits;
  reg [63:0] _RAND_4;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_5;
  reg  outputLengthCommitted;
  reg [31:0] _RAND_6;
  reg [63:0] inputMemAddr;
  reg [63:0] _RAND_7;
  reg [63:0] outputMemAddr;
  reg [63:0] _RAND_8;
  reg [63:0] outputLenAddr;
  reg [63:0] _RAND_9;
  reg  inputAddressAccepted;
  reg [31:0] _RAND_10;
  wire  _T_41;
  wire  _T_42;
  wire  _T_44;
  wire  _T_46;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_53;
  wire  _GEN_0;
  wire  inputBlockReadable;
  wire  _T_56;
  wire  _T_57;
  wire  _T_59;
  wire [9:0] _T_61;
  wire [9:0] _T_62;
  wire  _T_64;
  wire [47:0] _T_65;
  wire [63:0] _T_66;
  wire [63:0] _GEN_1;
  wire  _T_68;
  wire [31:0] _T_69;
  wire [47:0] _T_70;
  wire [15:0] _T_71;
  wire [63:0] _T_72;
  wire [63:0] _GEN_2;
  wire  _T_74;
  wire [15:0] _T_75;
  wire [31:0] _T_76;
  wire [31:0] _T_77;
  wire [63:0] _T_78;
  wire [63:0] _GEN_3;
  wire  _T_80;
  wire [47:0] _T_81;
  wire [63:0] _T_82;
  wire [63:0] _GEN_4;
  wire  _T_84;
  wire [47:0] _T_85;
  wire [63:0] _T_86;
  wire [63:0] _GEN_5;
  wire  _T_88;
  wire [31:0] _T_89;
  wire [47:0] _T_90;
  wire [15:0] _T_91;
  wire [63:0] _T_92;
  wire [63:0] _GEN_6;
  wire  _T_94;
  wire [15:0] _T_95;
  wire [31:0] _T_96;
  wire [31:0] _T_97;
  wire [63:0] _T_98;
  wire [63:0] _GEN_7;
  wire  _T_100;
  wire [47:0] _T_101;
  wire [63:0] _T_102;
  wire [63:0] _GEN_8;
  wire  _T_104;
  wire [47:0] _T_105;
  wire [63:0] _T_106;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire  _T_108;
  wire [31:0] _T_109;
  wire [47:0] _T_110;
  wire [15:0] _T_111;
  wire [63:0] _T_112;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire  _T_114;
  wire [15:0] _T_115;
  wire [31:0] _T_116;
  wire [31:0] _T_117;
  wire [63:0] _T_118;
  wire [63:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire  _T_120;
  wire [47:0] _T_121;
  wire [63:0] _T_122;
  wire [63:0] _GEN_15;
  wire [63:0] _GEN_16;
  wire  _T_124;
  wire [64:0] _T_128;
  wire [63:0] _T_129;
  wire  _GEN_17;
  wire  _GEN_18;
  wire [63:0] _GEN_19;
  wire [64:0] _T_135;
  wire [64:0] _T_136;
  wire [63:0] _T_137;
  wire [63:0] _T_139;
  wire [64:0] _T_141;
  wire [63:0] _T_142;
  wire [63:0] _GEN_20;
  wire [63:0] _GEN_21;
  wire [63:0] _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [63:0] _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire [63:0] _GEN_29;
  wire [63:0] _GEN_30;
  wire [63:0] _GEN_31;
  wire [63:0] _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _T_150;
  wire  _GEN_36;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_11;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_12;
  wire  _GEN_37;
  wire [63:0] _T_157;
  wire  _T_159;
  wire  _T_161;
  wire  _T_162;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _GEN_38;
  wire  _T_171;
  wire [4:0] _GEN_39;
  wire [5:0] _T_174;
  wire [4:0] _T_175;
  wire [4:0] _GEN_40;
  wire [4:0] _GEN_41;
  wire [15:0] outputBitsBlock;
  wire  _T_178;
  wire [15:0] _T_179;
  wire  _T_181;
  wire [15:0] _T_182;
  wire  _T_184;
  wire [15:0] _T_185;
  wire  _T_187;
  wire [15:0] _T_188;
  wire [15:0] _T_190;
  wire [15:0] _T_191;
  wire [15:0] _T_192;
  wire [15:0] _T_193;
  wire [15:0] _T_194;
  wire  _T_195;
  wire  _T_199;
  wire [63:0] _GEN_50;
  wire [64:0] _T_203;
  wire [63:0] _T_204;
  wire  _GEN_42;
  wire [63:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire [63:0] _GEN_48;
  wire [63:0] _GEN_49;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign _T_41 = inputAddressAccepted == 1'h0;
  assign _T_42 = initDone & core_io_inputMemConsumed;
  assign _T_44 = inputBitsRemaining == 64'h0;
  assign _T_46 = _T_44 == 1'h0;
  assign _T_47 = _T_42 & _T_46;
  assign _T_48 = isInit | _T_47;
  assign _T_49 = _T_41 & _T_48;
  assign _T_50 = io_inputMemAddrValid & io_inputMemAddrReady;
  assign _T_53 = reset == 1'h0;
  assign _GEN_0 = _T_50 ? 1'h1 : inputAddressAccepted;
  assign _T_56 = inputAddressAccepted & io_inputMemBlockValid;
  assign _T_57 = inputBlockReadable & initDone;
  assign _T_59 = inputBitsRemaining > 64'h200;
  assign _T_61 = inputBitsRemaining[9:0];
  assign _T_62 = _T_59 ? 10'h200 : _T_61;
  assign _T_64 = io_inputMemIdx == 5'h0;
  assign _T_65 = inputMemAddr[63:16];
  assign _T_66 = {_T_65,io_inputMemBlock};
  assign _GEN_1 = _T_64 ? _T_66 : inputMemAddr;
  assign _T_68 = io_inputMemIdx == 5'h1;
  assign _T_69 = inputMemAddr[63:32];
  assign _T_70 = {_T_69,io_inputMemBlock};
  assign _T_71 = inputMemAddr[15:0];
  assign _T_72 = {_T_70,_T_71};
  assign _GEN_2 = _T_68 ? _T_72 : _GEN_1;
  assign _T_74 = io_inputMemIdx == 5'h2;
  assign _T_75 = inputMemAddr[63:48];
  assign _T_76 = {_T_75,io_inputMemBlock};
  assign _T_77 = inputMemAddr[31:0];
  assign _T_78 = {_T_76,_T_77};
  assign _GEN_3 = _T_74 ? _T_78 : _GEN_2;
  assign _T_80 = io_inputMemIdx == 5'h3;
  assign _T_81 = inputMemAddr[47:0];
  assign _T_82 = {io_inputMemBlock,_T_81};
  assign _GEN_4 = _T_80 ? _T_82 : _GEN_3;
  assign _T_84 = io_inputMemIdx == 5'h4;
  assign _T_85 = inputBitsRemaining[63:16];
  assign _T_86 = {_T_85,io_inputMemBlock};
  assign _GEN_5 = _T_84 ? _T_86 : inputBitsRemaining;
  assign _T_88 = io_inputMemIdx == 5'h5;
  assign _T_89 = inputBitsRemaining[63:32];
  assign _T_90 = {_T_89,io_inputMemBlock};
  assign _T_91 = inputBitsRemaining[15:0];
  assign _T_92 = {_T_90,_T_91};
  assign _GEN_6 = _T_88 ? _T_92 : _GEN_5;
  assign _T_94 = io_inputMemIdx == 5'h6;
  assign _T_95 = inputBitsRemaining[63:48];
  assign _T_96 = {_T_95,io_inputMemBlock};
  assign _T_97 = inputBitsRemaining[31:0];
  assign _T_98 = {_T_96,_T_97};
  assign _GEN_7 = _T_94 ? _T_98 : _GEN_6;
  assign _T_100 = io_inputMemIdx == 5'h7;
  assign _T_101 = inputBitsRemaining[47:0];
  assign _T_102 = {io_inputMemBlock,_T_101};
  assign _GEN_8 = _T_100 ? _T_102 : _GEN_7;
  assign _T_104 = io_inputMemIdx == 5'h8;
  assign _T_105 = outputMemAddr[63:16];
  assign _T_106 = {_T_105,io_inputMemBlock};
  assign _GEN_9 = _T_104 ? _T_106 : outputMemAddr;
  assign _GEN_10 = _T_104 ? _T_106 : outputLenAddr;
  assign _T_108 = io_inputMemIdx == 5'h9;
  assign _T_109 = outputMemAddr[63:32];
  assign _T_110 = {_T_109,io_inputMemBlock};
  assign _T_111 = outputMemAddr[15:0];
  assign _T_112 = {_T_110,_T_111};
  assign _GEN_11 = _T_108 ? _T_112 : _GEN_9;
  assign _GEN_12 = _T_108 ? _T_112 : _GEN_10;
  assign _T_114 = io_inputMemIdx == 5'ha;
  assign _T_115 = outputMemAddr[63:48];
  assign _T_116 = {_T_115,io_inputMemBlock};
  assign _T_117 = outputMemAddr[31:0];
  assign _T_118 = {_T_116,_T_117};
  assign _GEN_13 = _T_114 ? _T_118 : _GEN_11;
  assign _GEN_14 = _T_114 ? _T_118 : _GEN_12;
  assign _T_120 = io_inputMemIdx == 5'hb;
  assign _T_121 = outputMemAddr[47:0];
  assign _T_122 = {io_inputMemBlock,_T_121};
  assign _GEN_15 = _T_120 ? _T_122 : _GEN_13;
  assign _GEN_16 = _T_120 ? _T_122 : _GEN_14;
  assign _T_124 = io_inputMemIdx == 5'h1f;
  assign _T_128 = outputMemAddr + 64'h40;
  assign _T_129 = _T_128[63:0];
  assign _GEN_17 = _T_124 ? 1'h0 : isInit;
  assign _GEN_18 = _T_124 ? 1'h1 : initDone;
  assign _GEN_19 = _T_124 ? _T_129 : _GEN_15;
  assign _T_135 = inputBitsRemaining - 64'h200;
  assign _T_136 = $unsigned(_T_135);
  assign _T_137 = _T_136[63:0];
  assign _T_139 = _T_59 ? _T_137 : 64'h0;
  assign _T_141 = inputMemAddr + 64'h40;
  assign _T_142 = _T_141[63:0];
  assign _GEN_20 = _T_124 ? _T_139 : inputBitsRemaining;
  assign _GEN_21 = _T_124 ? _T_142 : inputMemAddr;
  assign _GEN_22 = isInit ? _GEN_4 : _GEN_21;
  assign _GEN_23 = isInit ? _GEN_8 : _GEN_20;
  assign _GEN_24 = isInit ? _GEN_19 : outputMemAddr;
  assign _GEN_25 = isInit ? _GEN_16 : outputLenAddr;
  assign _GEN_26 = isInit ? _GEN_17 : isInit;
  assign _GEN_27 = isInit ? _GEN_18 : initDone;
  assign _GEN_28 = _T_124 ? 1'h0 : _GEN_0;
  assign _GEN_29 = inputBlockReadable ? _GEN_22 : inputMemAddr;
  assign _GEN_30 = inputBlockReadable ? _GEN_23 : inputBitsRemaining;
  assign _GEN_31 = inputBlockReadable ? _GEN_24 : outputMemAddr;
  assign _GEN_32 = inputBlockReadable ? _GEN_25 : outputLenAddr;
  assign _GEN_33 = inputBlockReadable ? _GEN_26 : isInit;
  assign _GEN_34 = inputBlockReadable ? _GEN_27 : initDone;
  assign _GEN_35 = inputBlockReadable ? _GEN_28 : _GEN_0;
  assign _T_150 = core_io_inputMemConsumed & _T_44;
  assign _GEN_36 = _T_150 ? 1'h1 : coreInputFinished;
  assign _GEN_37 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_157 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_159 = outputAddressAccepted == 1'h0;
  assign _T_161 = outputLengthCommitted == 1'h0;
  assign _T_162 = core_io_outputFinished & _T_161;
  assign _T_163 = core_io_outputMemBlockValid | _T_162;
  assign _T_164 = _T_159 & _T_163;
  assign _T_165 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_38 = _T_165 ? 1'h1 : outputAddressAccepted;
  assign _T_171 = outputBlockCounter == 5'h1f;
  assign _GEN_39 = io_outputMemBlockReady ? 5'h0 : outputBlockCounter;
  assign _T_174 = outputBlockCounter + 5'h1;
  assign _T_175 = _T_174[4:0];
  assign _GEN_40 = _T_171 ? _GEN_39 : _T_175;
  assign _GEN_41 = outputAddressAcceptedNext ? _GEN_40 : outputBlockCounter;
  assign _T_178 = outputBlockCounter == 5'h0;
  assign _T_179 = outputBits[15:0];
  assign _T_181 = outputBlockCounter == 5'h1;
  assign _T_182 = outputBits[31:16];
  assign _T_184 = outputBlockCounter == 5'h2;
  assign _T_185 = outputBits[47:32];
  assign _T_187 = outputBlockCounter == 5'h3;
  assign _T_188 = outputBits[63:48];
  assign _T_190 = _T_187 ? _T_188 : 16'h0;
  assign _T_191 = _T_184 ? _T_185 : _T_190;
  assign _T_192 = _T_181 ? _T_182 : _T_191;
  assign _T_193 = _T_178 ? _T_179 : _T_192;
  assign _T_194 = core_io_outputFinished ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_195 = outputAddressAcceptedNext & io_outputMemBlockReady;
  assign _T_199 = _T_195 & _T_171;
  assign _GEN_50 = {{54'd0}, core_io_outputBits};
  assign _T_203 = outputBits + _GEN_50;
  assign _T_204 = _T_203[63:0];
  assign _GEN_42 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _GEN_43 = core_io_outputFinished ? outputBits : _T_204;
  assign _GEN_44 = core_io_outputFinished ? _GEN_31 : _T_129;
  assign _GEN_45 = _T_199 ? 1'h0 : _GEN_38;
  assign _GEN_46 = _T_199 ? 1'h0 : _GEN_37;
  assign _GEN_47 = _T_199 ? _GEN_42 : outputLengthCommitted;
  assign _GEN_48 = _T_199 ? _GEN_43 : outputBits;
  assign _GEN_49 = _T_199 ? _GEN_44 : _GEN_31;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemAddrValid = _T_49;
  assign io_inputMemBlockReady = inputAddressAccepted;
  assign io_outputMemAddr = _T_157;
  assign io_outputMemAddrValid = _T_164;
  assign io_outputMemBlock = _T_194;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_inputFinished = _T_44;
  assign io_outputFinished = outputLengthCommitted;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_57;
  assign core_io_inputBits = _T_62;
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_io_outputMemFlushed = _T_195;
  assign core_clock = clock;
  assign core_reset = reset;
  assign inputBlockReadable = _T_56;
  assign outputBitsBlock = _T_193;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{$random}};
  inputBitsRemaining = _RAND_2[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  coreInputFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{$random}};
  outputBits = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputBlockCounter = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputLengthCommitted = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{$random}};
  inputMemAddr = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{$random}};
  outputMemAddr = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{$random}};
  outputLenAddr = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputAddressAccepted = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  outputAddressAccepted = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  outputAddressAcceptedNext = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 64'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_100) begin
            inputBitsRemaining <= _T_102;
          end else begin
            if (_T_94) begin
              inputBitsRemaining <= _T_98;
            end else begin
              if (_T_88) begin
                inputBitsRemaining <= _T_92;
              end else begin
                if (_T_84) begin
                  inputBitsRemaining <= _T_86;
                end
              end
            end
          end
        end else begin
          if (_T_124) begin
            if (_T_59) begin
              inputBitsRemaining <= _T_137;
            end else begin
              inputBitsRemaining <= 64'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_150) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 64'h0;
    end else begin
      if (_T_199) begin
        if (!(core_io_outputFinished)) begin
          outputBits <= _T_204;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_171) begin
          if (io_outputMemBlockReady) begin
            outputBlockCounter <= 5'h0;
          end
        end else begin
          outputBlockCounter <= _T_175;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_199) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 64'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_80) begin
            inputMemAddr <= _T_82;
          end else begin
            if (_T_74) begin
              inputMemAddr <= _T_78;
            end else begin
              if (_T_68) begin
                inputMemAddr <= _T_72;
              end else begin
                if (_T_64) begin
                  inputMemAddr <= _T_66;
                end
              end
            end
          end
        end else begin
          if (_T_124) begin
            inputMemAddr <= _T_142;
          end
        end
      end
    end
    if (_T_199) begin
      if (core_io_outputFinished) begin
        if (inputBlockReadable) begin
          if (isInit) begin
            if (_T_124) begin
              outputMemAddr <= _T_129;
            end else begin
              if (_T_120) begin
                outputMemAddr <= _T_122;
              end else begin
                if (_T_114) begin
                  outputMemAddr <= _T_118;
                end else begin
                  if (_T_108) begin
                    outputMemAddr <= _T_112;
                  end else begin
                    if (_T_104) begin
                      outputMemAddr <= _T_106;
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        outputMemAddr <= _T_129;
      end
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            outputMemAddr <= _T_129;
          end else begin
            if (_T_120) begin
              outputMemAddr <= _T_122;
            end else begin
              if (_T_114) begin
                outputMemAddr <= _T_118;
              end else begin
                if (_T_108) begin
                  outputMemAddr <= _T_112;
                end else begin
                  if (_T_104) begin
                    outputMemAddr <= _T_106;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (inputBlockReadable) begin
      if (isInit) begin
        if (_T_120) begin
          outputLenAddr <= _T_122;
        end else begin
          if (_T_114) begin
            outputLenAddr <= _T_118;
          end else begin
            if (_T_108) begin
              outputLenAddr <= _T_112;
            end else begin
              if (_T_104) begin
                outputLenAddr <= _T_106;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      inputAddressAccepted <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (_T_124) begin
          inputAddressAccepted <= 1'h0;
        end else begin
          if (_T_50) begin
            inputAddressAccepted <= 1'h1;
          end
        end
      end else begin
        if (_T_50) begin
          inputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_199) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_165) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_199) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_50 & _T_53) begin
          $fwrite(32'h80000002,"input address 0x%h accepted for core 1\n",io_inputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_165 & _T_53) begin
          $fwrite(32'h80000002,"output address 0x%h accepted for core 1\n",io_outputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module StreamingWrapper(
  input          clock,
  input          reset,
  output [63:0]  io_inputMemAddrs_0,
  output [63:0]  io_inputMemAddrs_1,
  output         io_inputMemAddrValids_0,
  output         io_inputMemAddrValids_1,
  input          io_inputMemAddrReadys_0,
  input          io_inputMemAddrReadys_1,
  input  [511:0] io_inputMemBlocks_0,
  input  [511:0] io_inputMemBlocks_1,
  input          io_inputMemBlockValids_0,
  input          io_inputMemBlockValids_1,
  output         io_inputMemBlockReadys_0,
  output         io_inputMemBlockReadys_1,
  output [63:0]  io_outputMemAddrs_0,
  output [63:0]  io_outputMemAddrs_1,
  output         io_outputMemAddrValids_0,
  output         io_outputMemAddrValids_1,
  input          io_outputMemAddrReadys_0,
  input          io_outputMemAddrReadys_1,
  output [511:0] io_outputMemBlocks_0,
  output [511:0] io_outputMemBlocks_1,
  output         io_outputMemBlockValids_0,
  output         io_outputMemBlockValids_1,
  input          io_outputMemBlockReadys_0,
  input          io_outputMemBlockReadys_1,
  output         io_finished
);
  wire  StreamingCore_clock;
  wire  StreamingCore_reset;
  wire [63:0] StreamingCore_io_inputMemAddr;
  wire  StreamingCore_io_inputMemAddrValid;
  wire  StreamingCore_io_inputMemAddrReady;
  wire [15:0] StreamingCore_io_inputMemBlock;
  wire [4:0] StreamingCore_io_inputMemIdx;
  wire  StreamingCore_io_inputMemBlockValid;
  wire  StreamingCore_io_inputMemBlockReady;
  wire [63:0] StreamingCore_io_outputMemAddr;
  wire  StreamingCore_io_outputMemAddrValid;
  wire  StreamingCore_io_outputMemAddrReady;
  wire [15:0] StreamingCore_io_outputMemBlock;
  wire [4:0] StreamingCore_io_outputMemIdx;
  wire  StreamingCore_io_outputMemBlockValid;
  wire  StreamingCore_io_outputMemBlockReady;
  wire  StreamingCore_io_inputFinished;
  wire  StreamingCore_io_outputFinished;
  wire  StreamingCore_1_clock;
  wire  StreamingCore_1_reset;
  wire [63:0] StreamingCore_1_io_inputMemAddr;
  wire  StreamingCore_1_io_inputMemAddrValid;
  wire  StreamingCore_1_io_inputMemAddrReady;
  wire [15:0] StreamingCore_1_io_inputMemBlock;
  wire [4:0] StreamingCore_1_io_inputMemIdx;
  wire  StreamingCore_1_io_inputMemBlockValid;
  wire  StreamingCore_1_io_inputMemBlockReady;
  wire [63:0] StreamingCore_1_io_outputMemAddr;
  wire  StreamingCore_1_io_outputMemAddrValid;
  wire  StreamingCore_1_io_outputMemAddrReady;
  wire [15:0] StreamingCore_1_io_outputMemBlock;
  wire [4:0] StreamingCore_1_io_outputMemIdx;
  wire  StreamingCore_1_io_outputMemBlockValid;
  wire  StreamingCore_1_io_outputMemBlockReady;
  wire  StreamingCore_1_io_inputFinished;
  wire  StreamingCore_1_io_outputFinished;
  wire [63:0] cores_0_inputMemAddr;
  wire  cores_0_inputMemAddrValid;
  wire  cores_0_inputMemAddrReady;
  wire [15:0] cores_0_inputMemBlock;
  wire [4:0] cores_0_inputMemIdx;
  wire  cores_0_inputMemBlockValid;
  wire  cores_0_inputMemBlockReady;
  wire [63:0] cores_0_outputMemAddr;
  wire  cores_0_outputMemAddrValid;
  wire  cores_0_outputMemAddrReady;
  wire [15:0] cores_0_outputMemBlock;
  wire [4:0] cores_0_outputMemIdx;
  wire  cores_0_outputMemBlockValid;
  wire  cores_0_outputMemBlockReady;
  wire  cores_0_inputFinished;
  wire  cores_0_outputFinished;
  wire [63:0] cores_1_inputMemAddr;
  wire  cores_1_inputMemAddrValid;
  wire  cores_1_inputMemAddrReady;
  wire [15:0] cores_1_inputMemBlock;
  wire [4:0] cores_1_inputMemIdx;
  wire  cores_1_inputMemBlockValid;
  wire  cores_1_inputMemBlockReady;
  wire [63:0] cores_1_outputMemAddr;
  wire  cores_1_outputMemAddrValid;
  wire  cores_1_outputMemAddrReady;
  wire [15:0] cores_1_outputMemBlock;
  wire [4:0] cores_1_outputMemIdx;
  wire  cores_1_outputMemBlockValid;
  wire  cores_1_outputMemBlockReady;
  wire  cores_1_inputFinished;
  wire  cores_1_outputFinished;
  reg [63:0] _T_238;
  reg [63:0] _RAND_0;
  reg  _T_240;
  reg [31:0] _RAND_1;
  reg  _T_242;
  reg [31:0] _RAND_2;
  reg  _T_244;
  reg [31:0] _RAND_3;
  reg [63:0] _T_246;
  reg [63:0] _RAND_4;
  reg  _T_248;
  reg [31:0] _RAND_5;
  reg  _T_250;
  reg [31:0] _RAND_6;
  reg  _T_252;
  reg [31:0] _RAND_7;
  reg [63:0] _T_254;
  reg [63:0] _RAND_8;
  reg  _T_256;
  reg [31:0] _RAND_9;
  reg  _T_258;
  reg [31:0] _RAND_10;
  reg [15:0] _T_260;
  reg [31:0] _RAND_11;
  reg [4:0] _T_262;
  reg [31:0] _RAND_12;
  reg  _T_264;
  reg [31:0] _RAND_13;
  reg [63:0] _T_266;
  reg [63:0] _RAND_14;
  reg  _T_268;
  reg [31:0] _RAND_15;
  reg  _T_270;
  reg [31:0] _RAND_16;
  reg [15:0] _T_272;
  reg [31:0] _RAND_17;
  reg [4:0] _T_274;
  reg [31:0] _RAND_18;
  reg  _T_276;
  reg [31:0] _RAND_19;
  reg  _T_279;
  reg [31:0] _RAND_20;
  reg  _T_282;
  reg [31:0] _RAND_21;
  reg  _T_285;
  reg [31:0] _RAND_22;
  reg  _T_288;
  reg [31:0] _RAND_23;
  reg  _T_291;
  reg [31:0] _RAND_24;
  wire  _T_293;
  wire [1:0] _T_295;
  wire  _T_296;
  wire  _GEN_4;
  reg  _T_299;
  reg [31:0] _RAND_25;
  reg  _T_302;
  reg [31:0] _RAND_26;
  reg [15:0] _T_306_0;
  reg [31:0] _RAND_27;
  reg [15:0] _T_306_1;
  reg [31:0] _RAND_28;
  reg [15:0] _T_306_2;
  reg [31:0] _RAND_29;
  reg [15:0] _T_306_3;
  reg [31:0] _RAND_30;
  reg [15:0] _T_306_4;
  reg [31:0] _RAND_31;
  reg [15:0] _T_306_5;
  reg [31:0] _RAND_32;
  reg [15:0] _T_306_6;
  reg [31:0] _RAND_33;
  reg [15:0] _T_306_7;
  reg [31:0] _RAND_34;
  reg [15:0] _T_306_8;
  reg [31:0] _RAND_35;
  reg [15:0] _T_306_9;
  reg [31:0] _RAND_36;
  reg [15:0] _T_306_10;
  reg [31:0] _RAND_37;
  reg [15:0] _T_306_11;
  reg [31:0] _RAND_38;
  reg [15:0] _T_306_12;
  reg [31:0] _RAND_39;
  reg [15:0] _T_306_13;
  reg [31:0] _RAND_40;
  reg [15:0] _T_306_14;
  reg [31:0] _RAND_41;
  reg [15:0] _T_306_15;
  reg [31:0] _RAND_42;
  reg [15:0] _T_306_16;
  reg [31:0] _RAND_43;
  reg [15:0] _T_306_17;
  reg [31:0] _RAND_44;
  reg [15:0] _T_306_18;
  reg [31:0] _RAND_45;
  reg [15:0] _T_306_19;
  reg [31:0] _RAND_46;
  reg [15:0] _T_306_20;
  reg [31:0] _RAND_47;
  reg [15:0] _T_306_21;
  reg [31:0] _RAND_48;
  reg [15:0] _T_306_22;
  reg [31:0] _RAND_49;
  reg [15:0] _T_306_23;
  reg [31:0] _RAND_50;
  reg [15:0] _T_306_24;
  reg [31:0] _RAND_51;
  reg [15:0] _T_306_25;
  reg [31:0] _RAND_52;
  reg [15:0] _T_306_26;
  reg [31:0] _RAND_53;
  reg [15:0] _T_306_27;
  reg [31:0] _RAND_54;
  reg [15:0] _T_306_28;
  reg [31:0] _RAND_55;
  reg [15:0] _T_306_29;
  reg [31:0] _RAND_56;
  reg [15:0] _T_306_30;
  reg [31:0] _RAND_57;
  reg [15:0] _T_306_31;
  reg [31:0] _RAND_58;
  reg [4:0] _T_343;
  reg [31:0] _RAND_59;
  reg  _T_346;
  reg [31:0] _RAND_60;
  wire  _T_347;
  wire [15:0] _T_348;
  wire [15:0] _T_349;
  wire [15:0] _T_350;
  wire [15:0] _T_351;
  wire [15:0] _T_352;
  wire [15:0] _T_353;
  wire [15:0] _T_354;
  wire [15:0] _T_355;
  wire [15:0] _T_356;
  wire [15:0] _T_357;
  wire [15:0] _T_358;
  wire [15:0] _T_359;
  wire [15:0] _T_360;
  wire [15:0] _T_361;
  wire [15:0] _T_362;
  wire [15:0] _T_363;
  wire [15:0] _T_364;
  wire [15:0] _T_365;
  wire [15:0] _T_366;
  wire [15:0] _T_367;
  wire [15:0] _T_368;
  wire [15:0] _T_369;
  wire [15:0] _T_370;
  wire [15:0] _T_371;
  wire [15:0] _T_372;
  wire [15:0] _T_373;
  wire [15:0] _T_374;
  wire [15:0] _T_375;
  wire [15:0] _T_376;
  wire [15:0] _T_377;
  wire [15:0] _T_378;
  wire [15:0] _T_379;
  wire  _T_383;
  wire [15:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire [15:0] _GEN_8;
  wire [15:0] _GEN_9;
  wire [15:0] _GEN_10;
  wire [15:0] _GEN_11;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_15;
  wire [15:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [15:0] _GEN_20;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_22;
  wire [15:0] _GEN_23;
  wire [15:0] _GEN_24;
  wire [15:0] _GEN_25;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  wire [15:0] _GEN_32;
  wire [15:0] _GEN_33;
  wire [15:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire [15:0] _GEN_36;
  wire  _GEN_37;
  wire  _T_385;
  wire [5:0] _T_389;
  wire [4:0] _T_390;
  wire  _GEN_38;
  wire [4:0] _GEN_39;
  wire  _GEN_40;
  wire [4:0] _GEN_41;
  wire  _T_393;
  wire  _T_395;
  wire  _T_396;
  wire  _GEN_42;
  wire  _T_398;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _T_403;
  wire  _T_405;
  wire  _T_407;
  wire [15:0] _GEN_0;
  wire [15:0] _GEN_45;
  wire [15:0] _GEN_46;
  wire [15:0] _GEN_47;
  wire [15:0] _GEN_48;
  wire [15:0] _GEN_49;
  wire [15:0] _GEN_50;
  wire [15:0] _GEN_51;
  wire [15:0] _GEN_52;
  wire [15:0] _GEN_53;
  wire [15:0] _GEN_54;
  wire [15:0] _GEN_55;
  wire [15:0] _GEN_56;
  wire [15:0] _GEN_57;
  wire [15:0] _GEN_58;
  wire [15:0] _GEN_59;
  wire [15:0] _GEN_60;
  wire [15:0] _GEN_61;
  wire [15:0] _GEN_62;
  wire [15:0] _GEN_63;
  wire [15:0] _GEN_64;
  wire [15:0] _GEN_65;
  wire [15:0] _GEN_66;
  wire [15:0] _GEN_67;
  wire [15:0] _GEN_68;
  wire [15:0] _GEN_69;
  wire [15:0] _GEN_70;
  wire [15:0] _GEN_71;
  wire [15:0] _GEN_72;
  wire [15:0] _GEN_73;
  wire [15:0] _GEN_74;
  wire [15:0] _GEN_75;
  wire  _T_412;
  wire  _T_417;
  wire  _T_418;
  wire [1:0] _T_423;
  wire  _T_424;
  wire  _T_425;
  wire  _GEN_76;
  wire  _GEN_77;
  wire  _GEN_78;
  reg  _T_430;
  reg [31:0] _RAND_61;
  wire  _T_432;
  wire [1:0] _T_434;
  wire  _T_435;
  wire  _GEN_79;
  reg  _T_438;
  reg [31:0] _RAND_62;
  reg  _T_441;
  reg [31:0] _RAND_63;
  reg [15:0] _T_445_0;
  reg [31:0] _RAND_64;
  reg [15:0] _T_445_1;
  reg [31:0] _RAND_65;
  reg [15:0] _T_445_2;
  reg [31:0] _RAND_66;
  reg [15:0] _T_445_3;
  reg [31:0] _RAND_67;
  reg [15:0] _T_445_4;
  reg [31:0] _RAND_68;
  reg [15:0] _T_445_5;
  reg [31:0] _RAND_69;
  reg [15:0] _T_445_6;
  reg [31:0] _RAND_70;
  reg [15:0] _T_445_7;
  reg [31:0] _RAND_71;
  reg [15:0] _T_445_8;
  reg [31:0] _RAND_72;
  reg [15:0] _T_445_9;
  reg [31:0] _RAND_73;
  reg [15:0] _T_445_10;
  reg [31:0] _RAND_74;
  reg [15:0] _T_445_11;
  reg [31:0] _RAND_75;
  reg [15:0] _T_445_12;
  reg [31:0] _RAND_76;
  reg [15:0] _T_445_13;
  reg [31:0] _RAND_77;
  reg [15:0] _T_445_14;
  reg [31:0] _RAND_78;
  reg [15:0] _T_445_15;
  reg [31:0] _RAND_79;
  reg [15:0] _T_445_16;
  reg [31:0] _RAND_80;
  reg [15:0] _T_445_17;
  reg [31:0] _RAND_81;
  reg [15:0] _T_445_18;
  reg [31:0] _RAND_82;
  reg [15:0] _T_445_19;
  reg [31:0] _RAND_83;
  reg [15:0] _T_445_20;
  reg [31:0] _RAND_84;
  reg [15:0] _T_445_21;
  reg [31:0] _RAND_85;
  reg [15:0] _T_445_22;
  reg [31:0] _RAND_86;
  reg [15:0] _T_445_23;
  reg [31:0] _RAND_87;
  reg [15:0] _T_445_24;
  reg [31:0] _RAND_88;
  reg [15:0] _T_445_25;
  reg [31:0] _RAND_89;
  reg [15:0] _T_445_26;
  reg [31:0] _RAND_90;
  reg [15:0] _T_445_27;
  reg [31:0] _RAND_91;
  reg [15:0] _T_445_28;
  reg [31:0] _RAND_92;
  reg [15:0] _T_445_29;
  reg [31:0] _RAND_93;
  reg [15:0] _T_445_30;
  reg [31:0] _RAND_94;
  reg [15:0] _T_445_31;
  reg [31:0] _RAND_95;
  reg [4:0] _T_482;
  reg [31:0] _RAND_96;
  reg  _T_485;
  reg [31:0] _RAND_97;
  wire  _T_486;
  wire [15:0] _T_487;
  wire [15:0] _T_488;
  wire [15:0] _T_489;
  wire [15:0] _T_490;
  wire [15:0] _T_491;
  wire [15:0] _T_492;
  wire [15:0] _T_493;
  wire [15:0] _T_494;
  wire [15:0] _T_495;
  wire [15:0] _T_496;
  wire [15:0] _T_497;
  wire [15:0] _T_498;
  wire [15:0] _T_499;
  wire [15:0] _T_500;
  wire [15:0] _T_501;
  wire [15:0] _T_502;
  wire [15:0] _T_503;
  wire [15:0] _T_504;
  wire [15:0] _T_505;
  wire [15:0] _T_506;
  wire [15:0] _T_507;
  wire [15:0] _T_508;
  wire [15:0] _T_509;
  wire [15:0] _T_510;
  wire [15:0] _T_511;
  wire [15:0] _T_512;
  wire [15:0] _T_513;
  wire [15:0] _T_514;
  wire [15:0] _T_515;
  wire [15:0] _T_516;
  wire [15:0] _T_517;
  wire [15:0] _T_518;
  wire [15:0] _GEN_80;
  wire [15:0] _GEN_81;
  wire [15:0] _GEN_82;
  wire [15:0] _GEN_83;
  wire [15:0] _GEN_84;
  wire [15:0] _GEN_85;
  wire [15:0] _GEN_86;
  wire [15:0] _GEN_87;
  wire [15:0] _GEN_88;
  wire [15:0] _GEN_89;
  wire [15:0] _GEN_90;
  wire [15:0] _GEN_91;
  wire [15:0] _GEN_92;
  wire [15:0] _GEN_93;
  wire [15:0] _GEN_94;
  wire [15:0] _GEN_95;
  wire [15:0] _GEN_96;
  wire [15:0] _GEN_97;
  wire [15:0] _GEN_98;
  wire [15:0] _GEN_99;
  wire [15:0] _GEN_100;
  wire [15:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire [15:0] _GEN_103;
  wire [15:0] _GEN_104;
  wire [15:0] _GEN_105;
  wire [15:0] _GEN_106;
  wire [15:0] _GEN_107;
  wire [15:0] _GEN_108;
  wire [15:0] _GEN_109;
  wire [15:0] _GEN_110;
  wire [15:0] _GEN_111;
  wire  _GEN_112;
  wire  _T_524;
  wire [5:0] _T_528;
  wire [4:0] _T_529;
  wire  _GEN_113;
  wire [4:0] _GEN_114;
  wire  _GEN_115;
  wire [4:0] _GEN_116;
  wire  _T_532;
  wire  _T_534;
  wire  _T_535;
  wire  _GEN_117;
  wire  _T_537;
  wire  _GEN_118;
  wire  _GEN_119;
  wire  _T_542;
  wire  _T_546;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_120;
  wire [15:0] _GEN_121;
  wire [15:0] _GEN_122;
  wire [15:0] _GEN_123;
  wire [15:0] _GEN_124;
  wire [15:0] _GEN_125;
  wire [15:0] _GEN_126;
  wire [15:0] _GEN_127;
  wire [15:0] _GEN_128;
  wire [15:0] _GEN_129;
  wire [15:0] _GEN_130;
  wire [15:0] _GEN_131;
  wire [15:0] _GEN_132;
  wire [15:0] _GEN_133;
  wire [15:0] _GEN_134;
  wire [15:0] _GEN_135;
  wire [15:0] _GEN_136;
  wire [15:0] _GEN_137;
  wire [15:0] _GEN_138;
  wire [15:0] _GEN_139;
  wire [15:0] _GEN_140;
  wire [15:0] _GEN_141;
  wire [15:0] _GEN_142;
  wire [15:0] _GEN_143;
  wire [15:0] _GEN_144;
  wire [15:0] _GEN_145;
  wire [15:0] _GEN_146;
  wire [15:0] _GEN_147;
  wire [15:0] _GEN_148;
  wire [15:0] _GEN_149;
  wire [15:0] _GEN_150;
  wire  _T_551;
  wire  _T_556;
  wire  _T_557;
  wire [1:0] _T_562;
  wire  _T_563;
  wire  _T_564;
  wire  _GEN_151;
  wire  _GEN_152;
  wire  _GEN_153;
  reg  _T_569;
  reg [31:0] _RAND_98;
  wire  _T_571;
  wire [1:0] _T_573;
  wire  _T_574;
  wire  _GEN_154;
  reg  _T_577;
  reg [31:0] _RAND_99;
  reg  _T_580;
  reg [31:0] _RAND_100;
  reg [15:0] _T_584_0;
  reg [31:0] _RAND_101;
  reg [15:0] _T_584_1;
  reg [31:0] _RAND_102;
  reg [15:0] _T_584_2;
  reg [31:0] _RAND_103;
  reg [15:0] _T_584_3;
  reg [31:0] _RAND_104;
  reg [15:0] _T_584_4;
  reg [31:0] _RAND_105;
  reg [15:0] _T_584_5;
  reg [31:0] _RAND_106;
  reg [15:0] _T_584_6;
  reg [31:0] _RAND_107;
  reg [15:0] _T_584_7;
  reg [31:0] _RAND_108;
  reg [15:0] _T_584_8;
  reg [31:0] _RAND_109;
  reg [15:0] _T_584_9;
  reg [31:0] _RAND_110;
  reg [15:0] _T_584_10;
  reg [31:0] _RAND_111;
  reg [15:0] _T_584_11;
  reg [31:0] _RAND_112;
  reg [15:0] _T_584_12;
  reg [31:0] _RAND_113;
  reg [15:0] _T_584_13;
  reg [31:0] _RAND_114;
  reg [15:0] _T_584_14;
  reg [31:0] _RAND_115;
  reg [15:0] _T_584_15;
  reg [31:0] _RAND_116;
  reg [15:0] _T_584_16;
  reg [31:0] _RAND_117;
  reg [15:0] _T_584_17;
  reg [31:0] _RAND_118;
  reg [15:0] _T_584_18;
  reg [31:0] _RAND_119;
  reg [15:0] _T_584_19;
  reg [31:0] _RAND_120;
  reg [15:0] _T_584_20;
  reg [31:0] _RAND_121;
  reg [15:0] _T_584_21;
  reg [31:0] _RAND_122;
  reg [15:0] _T_584_22;
  reg [31:0] _RAND_123;
  reg [15:0] _T_584_23;
  reg [31:0] _RAND_124;
  reg [15:0] _T_584_24;
  reg [31:0] _RAND_125;
  reg [15:0] _T_584_25;
  reg [31:0] _RAND_126;
  reg [15:0] _T_584_26;
  reg [31:0] _RAND_127;
  reg [15:0] _T_584_27;
  reg [31:0] _RAND_128;
  reg [15:0] _T_584_28;
  reg [31:0] _RAND_129;
  reg [15:0] _T_584_29;
  reg [31:0] _RAND_130;
  reg [15:0] _T_584_30;
  reg [31:0] _RAND_131;
  reg [15:0] _T_584_31;
  reg [31:0] _RAND_132;
  reg  _T_621;
  reg [31:0] _RAND_133;
  wire  _T_624;
  wire  _T_626;
  wire  _T_627;
  wire  _GEN_155;
  wire  _T_630;
  wire [15:0] _GEN_2;
  wire [15:0] _GEN_156;
  wire [15:0] _GEN_157;
  wire [15:0] _GEN_158;
  wire [15:0] _GEN_159;
  wire [15:0] _GEN_160;
  wire [15:0] _GEN_161;
  wire [15:0] _GEN_162;
  wire [15:0] _GEN_163;
  wire [15:0] _GEN_164;
  wire [15:0] _GEN_165;
  wire [15:0] _GEN_166;
  wire [15:0] _GEN_167;
  wire [15:0] _GEN_168;
  wire [15:0] _GEN_169;
  wire [15:0] _GEN_170;
  wire [15:0] _GEN_171;
  wire [15:0] _GEN_172;
  wire [15:0] _GEN_173;
  wire [15:0] _GEN_174;
  wire [15:0] _GEN_175;
  wire [15:0] _GEN_176;
  wire [15:0] _GEN_177;
  wire [15:0] _GEN_178;
  wire [15:0] _GEN_179;
  wire [15:0] _GEN_180;
  wire [15:0] _GEN_181;
  wire [15:0] _GEN_182;
  wire [15:0] _GEN_183;
  wire [15:0] _GEN_184;
  wire [15:0] _GEN_185;
  wire [15:0] _GEN_186;
  wire [15:0] _GEN_187;
  wire [15:0] _GEN_188;
  wire [15:0] _GEN_189;
  wire [15:0] _GEN_190;
  wire [15:0] _GEN_191;
  wire [15:0] _GEN_192;
  wire [15:0] _GEN_193;
  wire [15:0] _GEN_194;
  wire [15:0] _GEN_195;
  wire [15:0] _GEN_196;
  wire [15:0] _GEN_197;
  wire [15:0] _GEN_198;
  wire [15:0] _GEN_199;
  wire [15:0] _GEN_200;
  wire [15:0] _GEN_201;
  wire [15:0] _GEN_202;
  wire [15:0] _GEN_203;
  wire [15:0] _GEN_204;
  wire [15:0] _GEN_205;
  wire [15:0] _GEN_206;
  wire [15:0] _GEN_207;
  wire [15:0] _GEN_208;
  wire [15:0] _GEN_209;
  wire [15:0] _GEN_210;
  wire [15:0] _GEN_211;
  wire [15:0] _GEN_212;
  wire [15:0] _GEN_213;
  wire [15:0] _GEN_214;
  wire [15:0] _GEN_215;
  wire [15:0] _GEN_216;
  wire [15:0] _GEN_217;
  wire [15:0] _GEN_218;
  wire [15:0] _GEN_219;
  wire  _T_634;
  wire  _T_636;
  wire  _T_637;
  wire  _GEN_220;
  wire  _T_639;
  wire  _GEN_221;
  wire  _GEN_222;
  wire [31:0] _T_642;
  wire [31:0] _T_643;
  wire [63:0] _T_644;
  wire [31:0] _T_645;
  wire [31:0] _T_646;
  wire [63:0] _T_647;
  wire [127:0] _T_648;
  wire [31:0] _T_649;
  wire [31:0] _T_650;
  wire [63:0] _T_651;
  wire [31:0] _T_652;
  wire [31:0] _T_653;
  wire [63:0] _T_654;
  wire [127:0] _T_655;
  wire [255:0] _T_656;
  wire [31:0] _T_657;
  wire [31:0] _T_658;
  wire [63:0] _T_659;
  wire [31:0] _T_660;
  wire [31:0] _T_661;
  wire [63:0] _T_662;
  wire [127:0] _T_663;
  wire [31:0] _T_664;
  wire [31:0] _T_665;
  wire [63:0] _T_666;
  wire [31:0] _T_667;
  wire [31:0] _T_668;
  wire [63:0] _T_669;
  wire [127:0] _T_670;
  wire [255:0] _T_671;
  wire [511:0] _T_672;
  wire  _T_674;
  wire  _T_676;
  wire  _T_679;
  wire  _T_681;
  wire  _T_682;
  wire  _T_689;
  wire  _T_690;
  wire [1:0] _T_695;
  wire  _T_696;
  wire  _T_697;
  wire  _GEN_223;
  wire  _GEN_224;
  wire  _GEN_225;
  wire  _GEN_226;
  reg  _T_703;
  reg [31:0] _RAND_134;
  wire  _T_705;
  wire [1:0] _T_707;
  wire  _T_708;
  wire  _GEN_227;
  reg  _T_711;
  reg [31:0] _RAND_135;
  reg  _T_714;
  reg [31:0] _RAND_136;
  reg [15:0] _T_718_0;
  reg [31:0] _RAND_137;
  reg [15:0] _T_718_1;
  reg [31:0] _RAND_138;
  reg [15:0] _T_718_2;
  reg [31:0] _RAND_139;
  reg [15:0] _T_718_3;
  reg [31:0] _RAND_140;
  reg [15:0] _T_718_4;
  reg [31:0] _RAND_141;
  reg [15:0] _T_718_5;
  reg [31:0] _RAND_142;
  reg [15:0] _T_718_6;
  reg [31:0] _RAND_143;
  reg [15:0] _T_718_7;
  reg [31:0] _RAND_144;
  reg [15:0] _T_718_8;
  reg [31:0] _RAND_145;
  reg [15:0] _T_718_9;
  reg [31:0] _RAND_146;
  reg [15:0] _T_718_10;
  reg [31:0] _RAND_147;
  reg [15:0] _T_718_11;
  reg [31:0] _RAND_148;
  reg [15:0] _T_718_12;
  reg [31:0] _RAND_149;
  reg [15:0] _T_718_13;
  reg [31:0] _RAND_150;
  reg [15:0] _T_718_14;
  reg [31:0] _RAND_151;
  reg [15:0] _T_718_15;
  reg [31:0] _RAND_152;
  reg [15:0] _T_718_16;
  reg [31:0] _RAND_153;
  reg [15:0] _T_718_17;
  reg [31:0] _RAND_154;
  reg [15:0] _T_718_18;
  reg [31:0] _RAND_155;
  reg [15:0] _T_718_19;
  reg [31:0] _RAND_156;
  reg [15:0] _T_718_20;
  reg [31:0] _RAND_157;
  reg [15:0] _T_718_21;
  reg [31:0] _RAND_158;
  reg [15:0] _T_718_22;
  reg [31:0] _RAND_159;
  reg [15:0] _T_718_23;
  reg [31:0] _RAND_160;
  reg [15:0] _T_718_24;
  reg [31:0] _RAND_161;
  reg [15:0] _T_718_25;
  reg [31:0] _RAND_162;
  reg [15:0] _T_718_26;
  reg [31:0] _RAND_163;
  reg [15:0] _T_718_27;
  reg [31:0] _RAND_164;
  reg [15:0] _T_718_28;
  reg [31:0] _RAND_165;
  reg [15:0] _T_718_29;
  reg [31:0] _RAND_166;
  reg [15:0] _T_718_30;
  reg [31:0] _RAND_167;
  reg [15:0] _T_718_31;
  reg [31:0] _RAND_168;
  reg  _T_755;
  reg [31:0] _RAND_169;
  wire  _T_758;
  wire  _T_760;
  wire  _T_761;
  wire  _GEN_228;
  wire  _T_764;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_229;
  wire [15:0] _GEN_230;
  wire [15:0] _GEN_231;
  wire [15:0] _GEN_232;
  wire [15:0] _GEN_233;
  wire [15:0] _GEN_234;
  wire [15:0] _GEN_235;
  wire [15:0] _GEN_236;
  wire [15:0] _GEN_237;
  wire [15:0] _GEN_238;
  wire [15:0] _GEN_239;
  wire [15:0] _GEN_240;
  wire [15:0] _GEN_241;
  wire [15:0] _GEN_242;
  wire [15:0] _GEN_243;
  wire [15:0] _GEN_244;
  wire [15:0] _GEN_245;
  wire [15:0] _GEN_246;
  wire [15:0] _GEN_247;
  wire [15:0] _GEN_248;
  wire [15:0] _GEN_249;
  wire [15:0] _GEN_250;
  wire [15:0] _GEN_251;
  wire [15:0] _GEN_252;
  wire [15:0] _GEN_253;
  wire [15:0] _GEN_254;
  wire [15:0] _GEN_255;
  wire [15:0] _GEN_256;
  wire [15:0] _GEN_257;
  wire [15:0] _GEN_258;
  wire [15:0] _GEN_259;
  wire [15:0] _GEN_260;
  wire [15:0] _GEN_261;
  wire [15:0] _GEN_262;
  wire [15:0] _GEN_263;
  wire [15:0] _GEN_264;
  wire [15:0] _GEN_265;
  wire [15:0] _GEN_266;
  wire [15:0] _GEN_267;
  wire [15:0] _GEN_268;
  wire [15:0] _GEN_269;
  wire [15:0] _GEN_270;
  wire [15:0] _GEN_271;
  wire [15:0] _GEN_272;
  wire [15:0] _GEN_273;
  wire [15:0] _GEN_274;
  wire [15:0] _GEN_275;
  wire [15:0] _GEN_276;
  wire [15:0] _GEN_277;
  wire [15:0] _GEN_278;
  wire [15:0] _GEN_279;
  wire [15:0] _GEN_280;
  wire [15:0] _GEN_281;
  wire [15:0] _GEN_282;
  wire [15:0] _GEN_283;
  wire [15:0] _GEN_284;
  wire [15:0] _GEN_285;
  wire [15:0] _GEN_286;
  wire [15:0] _GEN_287;
  wire [15:0] _GEN_288;
  wire [15:0] _GEN_289;
  wire [15:0] _GEN_290;
  wire [15:0] _GEN_291;
  wire [15:0] _GEN_292;
  wire  _T_768;
  wire  _T_770;
  wire  _T_771;
  wire  _GEN_293;
  wire  _T_773;
  wire  _GEN_294;
  wire  _GEN_295;
  wire [31:0] _T_776;
  wire [31:0] _T_777;
  wire [63:0] _T_778;
  wire [31:0] _T_779;
  wire [31:0] _T_780;
  wire [63:0] _T_781;
  wire [127:0] _T_782;
  wire [31:0] _T_783;
  wire [31:0] _T_784;
  wire [63:0] _T_785;
  wire [31:0] _T_786;
  wire [31:0] _T_787;
  wire [63:0] _T_788;
  wire [127:0] _T_789;
  wire [255:0] _T_790;
  wire [31:0] _T_791;
  wire [31:0] _T_792;
  wire [63:0] _T_793;
  wire [31:0] _T_794;
  wire [31:0] _T_795;
  wire [63:0] _T_796;
  wire [127:0] _T_797;
  wire [31:0] _T_798;
  wire [31:0] _T_799;
  wire [63:0] _T_800;
  wire [31:0] _T_801;
  wire [31:0] _T_802;
  wire [63:0] _T_803;
  wire [127:0] _T_804;
  wire [255:0] _T_805;
  wire [511:0] _T_806;
  wire  _T_810;
  wire  _T_813;
  wire  _T_815;
  wire  _T_816;
  wire  _T_823;
  wire  _T_824;
  wire [1:0] _T_829;
  wire  _T_830;
  wire  _T_831;
  wire  _GEN_296;
  wire  _GEN_297;
  wire  _GEN_298;
  wire  _GEN_299;
  wire  cumFinished;
  StreamingCore StreamingCore (
    .clock(StreamingCore_clock),
    .reset(StreamingCore_reset),
    .io_inputMemAddr(StreamingCore_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_io_inputMemAddrValid),
    .io_inputMemAddrReady(StreamingCore_io_inputMemAddrReady),
    .io_inputMemBlock(StreamingCore_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_io_outputMemBlockReady),
    .io_inputFinished(StreamingCore_io_inputFinished),
    .io_outputFinished(StreamingCore_io_outputFinished)
  );
  StreamingCore_1 StreamingCore_1 (
    .clock(StreamingCore_1_clock),
    .reset(StreamingCore_1_reset),
    .io_inputMemAddr(StreamingCore_1_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_1_io_inputMemAddrValid),
    .io_inputMemAddrReady(StreamingCore_1_io_inputMemAddrReady),
    .io_inputMemBlock(StreamingCore_1_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_1_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_1_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_1_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_1_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_1_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_1_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_1_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_1_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_1_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_1_io_outputMemBlockReady),
    .io_inputFinished(StreamingCore_1_io_inputFinished),
    .io_outputFinished(StreamingCore_1_io_outputFinished)
  );
  assign _T_293 = _T_291 != 1'h1;
  assign _T_295 = _T_291 + 1'h1;
  assign _T_296 = _T_295[0:0];
  assign _GEN_4 = _T_293 ? _T_296 : _T_291;
  assign _T_347 = io_inputMemBlockReadys_0 & io_inputMemBlockValids_0;
  assign _T_348 = io_inputMemBlocks_0[15:0];
  assign _T_349 = io_inputMemBlocks_0[31:16];
  assign _T_350 = io_inputMemBlocks_0[47:32];
  assign _T_351 = io_inputMemBlocks_0[63:48];
  assign _T_352 = io_inputMemBlocks_0[79:64];
  assign _T_353 = io_inputMemBlocks_0[95:80];
  assign _T_354 = io_inputMemBlocks_0[111:96];
  assign _T_355 = io_inputMemBlocks_0[127:112];
  assign _T_356 = io_inputMemBlocks_0[143:128];
  assign _T_357 = io_inputMemBlocks_0[159:144];
  assign _T_358 = io_inputMemBlocks_0[175:160];
  assign _T_359 = io_inputMemBlocks_0[191:176];
  assign _T_360 = io_inputMemBlocks_0[207:192];
  assign _T_361 = io_inputMemBlocks_0[223:208];
  assign _T_362 = io_inputMemBlocks_0[239:224];
  assign _T_363 = io_inputMemBlocks_0[255:240];
  assign _T_364 = io_inputMemBlocks_0[271:256];
  assign _T_365 = io_inputMemBlocks_0[287:272];
  assign _T_366 = io_inputMemBlocks_0[303:288];
  assign _T_367 = io_inputMemBlocks_0[319:304];
  assign _T_368 = io_inputMemBlocks_0[335:320];
  assign _T_369 = io_inputMemBlocks_0[351:336];
  assign _T_370 = io_inputMemBlocks_0[367:352];
  assign _T_371 = io_inputMemBlocks_0[383:368];
  assign _T_372 = io_inputMemBlocks_0[399:384];
  assign _T_373 = io_inputMemBlocks_0[415:400];
  assign _T_374 = io_inputMemBlocks_0[431:416];
  assign _T_375 = io_inputMemBlocks_0[447:432];
  assign _T_376 = io_inputMemBlocks_0[463:448];
  assign _T_377 = io_inputMemBlocks_0[479:464];
  assign _T_378 = io_inputMemBlocks_0[495:480];
  assign _T_379 = io_inputMemBlocks_0[511:496];
  assign _T_383 = reset == 1'h0;
  assign _GEN_5 = _T_347 ? _T_348 : _T_306_0;
  assign _GEN_6 = _T_347 ? _T_349 : _T_306_1;
  assign _GEN_7 = _T_347 ? _T_350 : _T_306_2;
  assign _GEN_8 = _T_347 ? _T_351 : _T_306_3;
  assign _GEN_9 = _T_347 ? _T_352 : _T_306_4;
  assign _GEN_10 = _T_347 ? _T_353 : _T_306_5;
  assign _GEN_11 = _T_347 ? _T_354 : _T_306_6;
  assign _GEN_12 = _T_347 ? _T_355 : _T_306_7;
  assign _GEN_13 = _T_347 ? _T_356 : _T_306_8;
  assign _GEN_14 = _T_347 ? _T_357 : _T_306_9;
  assign _GEN_15 = _T_347 ? _T_358 : _T_306_10;
  assign _GEN_16 = _T_347 ? _T_359 : _T_306_11;
  assign _GEN_17 = _T_347 ? _T_360 : _T_306_12;
  assign _GEN_18 = _T_347 ? _T_361 : _T_306_13;
  assign _GEN_19 = _T_347 ? _T_362 : _T_306_14;
  assign _GEN_20 = _T_347 ? _T_363 : _T_306_15;
  assign _GEN_21 = _T_347 ? _T_364 : _T_306_16;
  assign _GEN_22 = _T_347 ? _T_365 : _T_306_17;
  assign _GEN_23 = _T_347 ? _T_366 : _T_306_18;
  assign _GEN_24 = _T_347 ? _T_367 : _T_306_19;
  assign _GEN_25 = _T_347 ? _T_368 : _T_306_20;
  assign _GEN_26 = _T_347 ? _T_369 : _T_306_21;
  assign _GEN_27 = _T_347 ? _T_370 : _T_306_22;
  assign _GEN_28 = _T_347 ? _T_371 : _T_306_23;
  assign _GEN_29 = _T_347 ? _T_372 : _T_306_24;
  assign _GEN_30 = _T_347 ? _T_373 : _T_306_25;
  assign _GEN_31 = _T_347 ? _T_374 : _T_306_26;
  assign _GEN_32 = _T_347 ? _T_375 : _T_306_27;
  assign _GEN_33 = _T_347 ? _T_376 : _T_306_28;
  assign _GEN_34 = _T_347 ? _T_377 : _T_306_29;
  assign _GEN_35 = _T_347 ? _T_378 : _T_306_30;
  assign _GEN_36 = _T_347 ? _T_379 : _T_306_31;
  assign _GEN_37 = _T_347 ? 1'h1 : _T_346;
  assign _T_385 = _T_343 == 5'h1f;
  assign _T_389 = _T_343 + 5'h1;
  assign _T_390 = _T_389[4:0];
  assign _GEN_38 = _T_385 ? 1'h0 : _GEN_37;
  assign _GEN_39 = _T_385 ? 5'h0 : _T_390;
  assign _GEN_40 = _T_346 ? _GEN_38 : _GEN_37;
  assign _GEN_41 = _T_346 ? _GEN_39 : _T_343;
  assign _T_393 = _T_291 & _T_240;
  assign _T_395 = _T_302 == 1'h0;
  assign _T_396 = _T_393 & _T_395;
  assign _GEN_42 = _T_396 ? 1'h1 : _T_299;
  assign _T_398 = _T_299 & io_inputMemAddrReadys_0;
  assign _GEN_43 = _T_398 ? 1'h0 : _GEN_42;
  assign _GEN_44 = _T_398 ? 1'h1 : _T_302;
  assign _T_403 = _T_291 & _T_242;
  assign _T_405 = _T_279 == 1'h0;
  assign _T_407 = _T_405 ? io_inputMemAddrReadys_0 : 1'h0;
  assign _GEN_45 = 5'h1 == _T_343 ? _T_306_1 : _T_306_0;
  assign _GEN_46 = 5'h2 == _T_343 ? _T_306_2 : _GEN_45;
  assign _GEN_47 = 5'h3 == _T_343 ? _T_306_3 : _GEN_46;
  assign _GEN_48 = 5'h4 == _T_343 ? _T_306_4 : _GEN_47;
  assign _GEN_49 = 5'h5 == _T_343 ? _T_306_5 : _GEN_48;
  assign _GEN_50 = 5'h6 == _T_343 ? _T_306_6 : _GEN_49;
  assign _GEN_51 = 5'h7 == _T_343 ? _T_306_7 : _GEN_50;
  assign _GEN_52 = 5'h8 == _T_343 ? _T_306_8 : _GEN_51;
  assign _GEN_53 = 5'h9 == _T_343 ? _T_306_9 : _GEN_52;
  assign _GEN_54 = 5'ha == _T_343 ? _T_306_10 : _GEN_53;
  assign _GEN_55 = 5'hb == _T_343 ? _T_306_11 : _GEN_54;
  assign _GEN_56 = 5'hc == _T_343 ? _T_306_12 : _GEN_55;
  assign _GEN_57 = 5'hd == _T_343 ? _T_306_13 : _GEN_56;
  assign _GEN_58 = 5'he == _T_343 ? _T_306_14 : _GEN_57;
  assign _GEN_59 = 5'hf == _T_343 ? _T_306_15 : _GEN_58;
  assign _GEN_60 = 5'h10 == _T_343 ? _T_306_16 : _GEN_59;
  assign _GEN_61 = 5'h11 == _T_343 ? _T_306_17 : _GEN_60;
  assign _GEN_62 = 5'h12 == _T_343 ? _T_306_18 : _GEN_61;
  assign _GEN_63 = 5'h13 == _T_343 ? _T_306_19 : _GEN_62;
  assign _GEN_64 = 5'h14 == _T_343 ? _T_306_20 : _GEN_63;
  assign _GEN_65 = 5'h15 == _T_343 ? _T_306_21 : _GEN_64;
  assign _GEN_66 = 5'h16 == _T_343 ? _T_306_22 : _GEN_65;
  assign _GEN_67 = 5'h17 == _T_343 ? _T_306_23 : _GEN_66;
  assign _GEN_68 = 5'h18 == _T_343 ? _T_306_24 : _GEN_67;
  assign _GEN_69 = 5'h19 == _T_343 ? _T_306_25 : _GEN_68;
  assign _GEN_70 = 5'h1a == _T_343 ? _T_306_26 : _GEN_69;
  assign _GEN_71 = 5'h1b == _T_343 ? _T_306_27 : _GEN_70;
  assign _GEN_72 = 5'h1c == _T_343 ? _T_306_28 : _GEN_71;
  assign _GEN_73 = 5'h1d == _T_343 ? _T_306_29 : _GEN_72;
  assign _GEN_74 = 5'h1e == _T_343 ? _T_306_30 : _GEN_73;
  assign _GEN_75 = 5'h1f == _T_343 ? _T_306_31 : _GEN_74;
  assign _T_412 = _T_405 ? _T_346 : 1'h0;
  assign _T_417 = _T_244 | _T_385;
  assign _T_418 = _T_291 & _T_417;
  assign _T_423 = _T_279 + 1'h1;
  assign _T_424 = _T_423[0:0];
  assign _T_425 = _T_405 ? 1'h0 : _T_424;
  assign _GEN_76 = _T_418 ? _T_425 : _T_279;
  assign _GEN_77 = _T_418 ? 1'h0 : _GEN_4;
  assign _GEN_78 = _T_418 ? 1'h0 : _GEN_44;
  assign _T_432 = _T_430 != 1'h1;
  assign _T_434 = _T_430 + 1'h1;
  assign _T_435 = _T_434[0:0];
  assign _GEN_79 = _T_432 ? _T_435 : _T_430;
  assign _T_486 = io_inputMemBlockReadys_1 & io_inputMemBlockValids_1;
  assign _T_487 = io_inputMemBlocks_1[15:0];
  assign _T_488 = io_inputMemBlocks_1[31:16];
  assign _T_489 = io_inputMemBlocks_1[47:32];
  assign _T_490 = io_inputMemBlocks_1[63:48];
  assign _T_491 = io_inputMemBlocks_1[79:64];
  assign _T_492 = io_inputMemBlocks_1[95:80];
  assign _T_493 = io_inputMemBlocks_1[111:96];
  assign _T_494 = io_inputMemBlocks_1[127:112];
  assign _T_495 = io_inputMemBlocks_1[143:128];
  assign _T_496 = io_inputMemBlocks_1[159:144];
  assign _T_497 = io_inputMemBlocks_1[175:160];
  assign _T_498 = io_inputMemBlocks_1[191:176];
  assign _T_499 = io_inputMemBlocks_1[207:192];
  assign _T_500 = io_inputMemBlocks_1[223:208];
  assign _T_501 = io_inputMemBlocks_1[239:224];
  assign _T_502 = io_inputMemBlocks_1[255:240];
  assign _T_503 = io_inputMemBlocks_1[271:256];
  assign _T_504 = io_inputMemBlocks_1[287:272];
  assign _T_505 = io_inputMemBlocks_1[303:288];
  assign _T_506 = io_inputMemBlocks_1[319:304];
  assign _T_507 = io_inputMemBlocks_1[335:320];
  assign _T_508 = io_inputMemBlocks_1[351:336];
  assign _T_509 = io_inputMemBlocks_1[367:352];
  assign _T_510 = io_inputMemBlocks_1[383:368];
  assign _T_511 = io_inputMemBlocks_1[399:384];
  assign _T_512 = io_inputMemBlocks_1[415:400];
  assign _T_513 = io_inputMemBlocks_1[431:416];
  assign _T_514 = io_inputMemBlocks_1[447:432];
  assign _T_515 = io_inputMemBlocks_1[463:448];
  assign _T_516 = io_inputMemBlocks_1[479:464];
  assign _T_517 = io_inputMemBlocks_1[495:480];
  assign _T_518 = io_inputMemBlocks_1[511:496];
  assign _GEN_80 = _T_486 ? _T_487 : _T_445_0;
  assign _GEN_81 = _T_486 ? _T_488 : _T_445_1;
  assign _GEN_82 = _T_486 ? _T_489 : _T_445_2;
  assign _GEN_83 = _T_486 ? _T_490 : _T_445_3;
  assign _GEN_84 = _T_486 ? _T_491 : _T_445_4;
  assign _GEN_85 = _T_486 ? _T_492 : _T_445_5;
  assign _GEN_86 = _T_486 ? _T_493 : _T_445_6;
  assign _GEN_87 = _T_486 ? _T_494 : _T_445_7;
  assign _GEN_88 = _T_486 ? _T_495 : _T_445_8;
  assign _GEN_89 = _T_486 ? _T_496 : _T_445_9;
  assign _GEN_90 = _T_486 ? _T_497 : _T_445_10;
  assign _GEN_91 = _T_486 ? _T_498 : _T_445_11;
  assign _GEN_92 = _T_486 ? _T_499 : _T_445_12;
  assign _GEN_93 = _T_486 ? _T_500 : _T_445_13;
  assign _GEN_94 = _T_486 ? _T_501 : _T_445_14;
  assign _GEN_95 = _T_486 ? _T_502 : _T_445_15;
  assign _GEN_96 = _T_486 ? _T_503 : _T_445_16;
  assign _GEN_97 = _T_486 ? _T_504 : _T_445_17;
  assign _GEN_98 = _T_486 ? _T_505 : _T_445_18;
  assign _GEN_99 = _T_486 ? _T_506 : _T_445_19;
  assign _GEN_100 = _T_486 ? _T_507 : _T_445_20;
  assign _GEN_101 = _T_486 ? _T_508 : _T_445_21;
  assign _GEN_102 = _T_486 ? _T_509 : _T_445_22;
  assign _GEN_103 = _T_486 ? _T_510 : _T_445_23;
  assign _GEN_104 = _T_486 ? _T_511 : _T_445_24;
  assign _GEN_105 = _T_486 ? _T_512 : _T_445_25;
  assign _GEN_106 = _T_486 ? _T_513 : _T_445_26;
  assign _GEN_107 = _T_486 ? _T_514 : _T_445_27;
  assign _GEN_108 = _T_486 ? _T_515 : _T_445_28;
  assign _GEN_109 = _T_486 ? _T_516 : _T_445_29;
  assign _GEN_110 = _T_486 ? _T_517 : _T_445_30;
  assign _GEN_111 = _T_486 ? _T_518 : _T_445_31;
  assign _GEN_112 = _T_486 ? 1'h1 : _T_485;
  assign _T_524 = _T_482 == 5'h1f;
  assign _T_528 = _T_482 + 5'h1;
  assign _T_529 = _T_528[4:0];
  assign _GEN_113 = _T_524 ? 1'h0 : _GEN_112;
  assign _GEN_114 = _T_524 ? 5'h0 : _T_529;
  assign _GEN_115 = _T_485 ? _GEN_113 : _GEN_112;
  assign _GEN_116 = _T_485 ? _GEN_114 : _T_482;
  assign _T_532 = _T_430 & _T_248;
  assign _T_534 = _T_441 == 1'h0;
  assign _T_535 = _T_532 & _T_534;
  assign _GEN_117 = _T_535 ? 1'h1 : _T_438;
  assign _T_537 = _T_438 & io_inputMemAddrReadys_1;
  assign _GEN_118 = _T_537 ? 1'h0 : _GEN_117;
  assign _GEN_119 = _T_537 ? 1'h1 : _T_441;
  assign _T_542 = _T_430 & _T_250;
  assign _T_546 = _T_282 ? io_inputMemAddrReadys_1 : 1'h0;
  assign _GEN_120 = 5'h1 == _T_482 ? _T_445_1 : _T_445_0;
  assign _GEN_121 = 5'h2 == _T_482 ? _T_445_2 : _GEN_120;
  assign _GEN_122 = 5'h3 == _T_482 ? _T_445_3 : _GEN_121;
  assign _GEN_123 = 5'h4 == _T_482 ? _T_445_4 : _GEN_122;
  assign _GEN_124 = 5'h5 == _T_482 ? _T_445_5 : _GEN_123;
  assign _GEN_125 = 5'h6 == _T_482 ? _T_445_6 : _GEN_124;
  assign _GEN_126 = 5'h7 == _T_482 ? _T_445_7 : _GEN_125;
  assign _GEN_127 = 5'h8 == _T_482 ? _T_445_8 : _GEN_126;
  assign _GEN_128 = 5'h9 == _T_482 ? _T_445_9 : _GEN_127;
  assign _GEN_129 = 5'ha == _T_482 ? _T_445_10 : _GEN_128;
  assign _GEN_130 = 5'hb == _T_482 ? _T_445_11 : _GEN_129;
  assign _GEN_131 = 5'hc == _T_482 ? _T_445_12 : _GEN_130;
  assign _GEN_132 = 5'hd == _T_482 ? _T_445_13 : _GEN_131;
  assign _GEN_133 = 5'he == _T_482 ? _T_445_14 : _GEN_132;
  assign _GEN_134 = 5'hf == _T_482 ? _T_445_15 : _GEN_133;
  assign _GEN_135 = 5'h10 == _T_482 ? _T_445_16 : _GEN_134;
  assign _GEN_136 = 5'h11 == _T_482 ? _T_445_17 : _GEN_135;
  assign _GEN_137 = 5'h12 == _T_482 ? _T_445_18 : _GEN_136;
  assign _GEN_138 = 5'h13 == _T_482 ? _T_445_19 : _GEN_137;
  assign _GEN_139 = 5'h14 == _T_482 ? _T_445_20 : _GEN_138;
  assign _GEN_140 = 5'h15 == _T_482 ? _T_445_21 : _GEN_139;
  assign _GEN_141 = 5'h16 == _T_482 ? _T_445_22 : _GEN_140;
  assign _GEN_142 = 5'h17 == _T_482 ? _T_445_23 : _GEN_141;
  assign _GEN_143 = 5'h18 == _T_482 ? _T_445_24 : _GEN_142;
  assign _GEN_144 = 5'h19 == _T_482 ? _T_445_25 : _GEN_143;
  assign _GEN_145 = 5'h1a == _T_482 ? _T_445_26 : _GEN_144;
  assign _GEN_146 = 5'h1b == _T_482 ? _T_445_27 : _GEN_145;
  assign _GEN_147 = 5'h1c == _T_482 ? _T_445_28 : _GEN_146;
  assign _GEN_148 = 5'h1d == _T_482 ? _T_445_29 : _GEN_147;
  assign _GEN_149 = 5'h1e == _T_482 ? _T_445_30 : _GEN_148;
  assign _GEN_150 = 5'h1f == _T_482 ? _T_445_31 : _GEN_149;
  assign _T_551 = _T_282 ? _T_485 : 1'h0;
  assign _T_556 = _T_252 | _T_524;
  assign _T_557 = _T_430 & _T_556;
  assign _T_562 = _T_282 + 1'h1;
  assign _T_563 = _T_562[0:0];
  assign _T_564 = _T_282 ? 1'h1 : _T_563;
  assign _GEN_151 = _T_557 ? _T_564 : _T_282;
  assign _GEN_152 = _T_557 ? 1'h0 : _GEN_79;
  assign _GEN_153 = _T_557 ? 1'h0 : _GEN_119;
  assign _T_571 = _T_569 != 1'h1;
  assign _T_573 = _T_569 + 1'h1;
  assign _T_574 = _T_573[0:0];
  assign _GEN_154 = _T_571 ? _T_574 : _T_569;
  assign _T_624 = _T_569 & _T_258;
  assign _T_626 = _T_262 == 5'h1f;
  assign _T_627 = _T_624 & _T_626;
  assign _GEN_155 = _T_627 ? 1'h1 : _T_621;
  assign _T_630 = _T_621 == 1'h0;
  assign _GEN_156 = 5'h0 == _T_262 ? _GEN_2 : _T_584_0;
  assign _GEN_157 = 5'h1 == _T_262 ? _GEN_2 : _T_584_1;
  assign _GEN_158 = 5'h2 == _T_262 ? _GEN_2 : _T_584_2;
  assign _GEN_159 = 5'h3 == _T_262 ? _GEN_2 : _T_584_3;
  assign _GEN_160 = 5'h4 == _T_262 ? _GEN_2 : _T_584_4;
  assign _GEN_161 = 5'h5 == _T_262 ? _GEN_2 : _T_584_5;
  assign _GEN_162 = 5'h6 == _T_262 ? _GEN_2 : _T_584_6;
  assign _GEN_163 = 5'h7 == _T_262 ? _GEN_2 : _T_584_7;
  assign _GEN_164 = 5'h8 == _T_262 ? _GEN_2 : _T_584_8;
  assign _GEN_165 = 5'h9 == _T_262 ? _GEN_2 : _T_584_9;
  assign _GEN_166 = 5'ha == _T_262 ? _GEN_2 : _T_584_10;
  assign _GEN_167 = 5'hb == _T_262 ? _GEN_2 : _T_584_11;
  assign _GEN_168 = 5'hc == _T_262 ? _GEN_2 : _T_584_12;
  assign _GEN_169 = 5'hd == _T_262 ? _GEN_2 : _T_584_13;
  assign _GEN_170 = 5'he == _T_262 ? _GEN_2 : _T_584_14;
  assign _GEN_171 = 5'hf == _T_262 ? _GEN_2 : _T_584_15;
  assign _GEN_172 = 5'h10 == _T_262 ? _GEN_2 : _T_584_16;
  assign _GEN_173 = 5'h11 == _T_262 ? _GEN_2 : _T_584_17;
  assign _GEN_174 = 5'h12 == _T_262 ? _GEN_2 : _T_584_18;
  assign _GEN_175 = 5'h13 == _T_262 ? _GEN_2 : _T_584_19;
  assign _GEN_176 = 5'h14 == _T_262 ? _GEN_2 : _T_584_20;
  assign _GEN_177 = 5'h15 == _T_262 ? _GEN_2 : _T_584_21;
  assign _GEN_178 = 5'h16 == _T_262 ? _GEN_2 : _T_584_22;
  assign _GEN_179 = 5'h17 == _T_262 ? _GEN_2 : _T_584_23;
  assign _GEN_180 = 5'h18 == _T_262 ? _GEN_2 : _T_584_24;
  assign _GEN_181 = 5'h19 == _T_262 ? _GEN_2 : _T_584_25;
  assign _GEN_182 = 5'h1a == _T_262 ? _GEN_2 : _T_584_26;
  assign _GEN_183 = 5'h1b == _T_262 ? _GEN_2 : _T_584_27;
  assign _GEN_184 = 5'h1c == _T_262 ? _GEN_2 : _T_584_28;
  assign _GEN_185 = 5'h1d == _T_262 ? _GEN_2 : _T_584_29;
  assign _GEN_186 = 5'h1e == _T_262 ? _GEN_2 : _T_584_30;
  assign _GEN_187 = 5'h1f == _T_262 ? _GEN_2 : _T_584_31;
  assign _GEN_188 = _T_630 ? _GEN_156 : _T_584_0;
  assign _GEN_189 = _T_630 ? _GEN_157 : _T_584_1;
  assign _GEN_190 = _T_630 ? _GEN_158 : _T_584_2;
  assign _GEN_191 = _T_630 ? _GEN_159 : _T_584_3;
  assign _GEN_192 = _T_630 ? _GEN_160 : _T_584_4;
  assign _GEN_193 = _T_630 ? _GEN_161 : _T_584_5;
  assign _GEN_194 = _T_630 ? _GEN_162 : _T_584_6;
  assign _GEN_195 = _T_630 ? _GEN_163 : _T_584_7;
  assign _GEN_196 = _T_630 ? _GEN_164 : _T_584_8;
  assign _GEN_197 = _T_630 ? _GEN_165 : _T_584_9;
  assign _GEN_198 = _T_630 ? _GEN_166 : _T_584_10;
  assign _GEN_199 = _T_630 ? _GEN_167 : _T_584_11;
  assign _GEN_200 = _T_630 ? _GEN_168 : _T_584_12;
  assign _GEN_201 = _T_630 ? _GEN_169 : _T_584_13;
  assign _GEN_202 = _T_630 ? _GEN_170 : _T_584_14;
  assign _GEN_203 = _T_630 ? _GEN_171 : _T_584_15;
  assign _GEN_204 = _T_630 ? _GEN_172 : _T_584_16;
  assign _GEN_205 = _T_630 ? _GEN_173 : _T_584_17;
  assign _GEN_206 = _T_630 ? _GEN_174 : _T_584_18;
  assign _GEN_207 = _T_630 ? _GEN_175 : _T_584_19;
  assign _GEN_208 = _T_630 ? _GEN_176 : _T_584_20;
  assign _GEN_209 = _T_630 ? _GEN_177 : _T_584_21;
  assign _GEN_210 = _T_630 ? _GEN_178 : _T_584_22;
  assign _GEN_211 = _T_630 ? _GEN_179 : _T_584_23;
  assign _GEN_212 = _T_630 ? _GEN_180 : _T_584_24;
  assign _GEN_213 = _T_630 ? _GEN_181 : _T_584_25;
  assign _GEN_214 = _T_630 ? _GEN_182 : _T_584_26;
  assign _GEN_215 = _T_630 ? _GEN_183 : _T_584_27;
  assign _GEN_216 = _T_630 ? _GEN_184 : _T_584_28;
  assign _GEN_217 = _T_630 ? _GEN_185 : _T_584_29;
  assign _GEN_218 = _T_630 ? _GEN_186 : _T_584_30;
  assign _GEN_219 = _T_630 ? _GEN_187 : _T_584_31;
  assign _T_634 = _T_569 & _T_256;
  assign _T_636 = _T_580 == 1'h0;
  assign _T_637 = _T_634 & _T_636;
  assign _GEN_220 = _T_637 ? 1'h1 : _T_577;
  assign _T_639 = _T_577 & io_outputMemAddrReadys_0;
  assign _GEN_221 = _T_639 ? 1'h0 : _GEN_220;
  assign _GEN_222 = _T_639 ? 1'h1 : _T_580;
  assign _T_642 = {_T_584_1,_T_584_0};
  assign _T_643 = {_T_584_3,_T_584_2};
  assign _T_644 = {_T_643,_T_642};
  assign _T_645 = {_T_584_5,_T_584_4};
  assign _T_646 = {_T_584_7,_T_584_6};
  assign _T_647 = {_T_646,_T_645};
  assign _T_648 = {_T_647,_T_644};
  assign _T_649 = {_T_584_9,_T_584_8};
  assign _T_650 = {_T_584_11,_T_584_10};
  assign _T_651 = {_T_650,_T_649};
  assign _T_652 = {_T_584_13,_T_584_12};
  assign _T_653 = {_T_584_15,_T_584_14};
  assign _T_654 = {_T_653,_T_652};
  assign _T_655 = {_T_654,_T_651};
  assign _T_656 = {_T_655,_T_648};
  assign _T_657 = {_T_584_17,_T_584_16};
  assign _T_658 = {_T_584_19,_T_584_18};
  assign _T_659 = {_T_658,_T_657};
  assign _T_660 = {_T_584_21,_T_584_20};
  assign _T_661 = {_T_584_23,_T_584_22};
  assign _T_662 = {_T_661,_T_660};
  assign _T_663 = {_T_662,_T_659};
  assign _T_664 = {_T_584_25,_T_584_24};
  assign _T_665 = {_T_584_27,_T_584_26};
  assign _T_666 = {_T_665,_T_664};
  assign _T_667 = {_T_584_29,_T_584_28};
  assign _T_668 = {_T_584_31,_T_584_30};
  assign _T_669 = {_T_668,_T_667};
  assign _T_670 = {_T_669,_T_666};
  assign _T_671 = {_T_670,_T_663};
  assign _T_672 = {_T_671,_T_656};
  assign _T_674 = _T_285 == 1'h0;
  assign _T_676 = _T_674 ? io_outputMemAddrReadys_0 : 1'h0;
  assign _T_679 = io_outputMemBlockReadys_0 & _T_621;
  assign _T_681 = _T_674 ? _T_679 : 1'h0;
  assign _T_682 = io_outputMemBlockReadys_0 & io_outputMemBlockValids_0;
  assign _T_689 = _T_264 | _T_679;
  assign _T_690 = _T_569 & _T_689;
  assign _T_695 = _T_285 + 1'h1;
  assign _T_696 = _T_695[0:0];
  assign _T_697 = _T_674 ? 1'h0 : _T_696;
  assign _GEN_223 = _T_690 ? _T_697 : _T_285;
  assign _GEN_224 = _T_690 ? 1'h0 : _GEN_155;
  assign _GEN_225 = _T_690 ? 1'h0 : _GEN_154;
  assign _GEN_226 = _T_690 ? 1'h0 : _GEN_222;
  assign _T_705 = _T_703 != 1'h1;
  assign _T_707 = _T_703 + 1'h1;
  assign _T_708 = _T_707[0:0];
  assign _GEN_227 = _T_705 ? _T_708 : _T_703;
  assign _T_758 = _T_703 & _T_270;
  assign _T_760 = _T_274 == 5'h1f;
  assign _T_761 = _T_758 & _T_760;
  assign _GEN_228 = _T_761 ? 1'h1 : _T_755;
  assign _T_764 = _T_755 == 1'h0;
  assign _GEN_229 = 5'h0 == _T_274 ? _GEN_3 : _T_718_0;
  assign _GEN_230 = 5'h1 == _T_274 ? _GEN_3 : _T_718_1;
  assign _GEN_231 = 5'h2 == _T_274 ? _GEN_3 : _T_718_2;
  assign _GEN_232 = 5'h3 == _T_274 ? _GEN_3 : _T_718_3;
  assign _GEN_233 = 5'h4 == _T_274 ? _GEN_3 : _T_718_4;
  assign _GEN_234 = 5'h5 == _T_274 ? _GEN_3 : _T_718_5;
  assign _GEN_235 = 5'h6 == _T_274 ? _GEN_3 : _T_718_6;
  assign _GEN_236 = 5'h7 == _T_274 ? _GEN_3 : _T_718_7;
  assign _GEN_237 = 5'h8 == _T_274 ? _GEN_3 : _T_718_8;
  assign _GEN_238 = 5'h9 == _T_274 ? _GEN_3 : _T_718_9;
  assign _GEN_239 = 5'ha == _T_274 ? _GEN_3 : _T_718_10;
  assign _GEN_240 = 5'hb == _T_274 ? _GEN_3 : _T_718_11;
  assign _GEN_241 = 5'hc == _T_274 ? _GEN_3 : _T_718_12;
  assign _GEN_242 = 5'hd == _T_274 ? _GEN_3 : _T_718_13;
  assign _GEN_243 = 5'he == _T_274 ? _GEN_3 : _T_718_14;
  assign _GEN_244 = 5'hf == _T_274 ? _GEN_3 : _T_718_15;
  assign _GEN_245 = 5'h10 == _T_274 ? _GEN_3 : _T_718_16;
  assign _GEN_246 = 5'h11 == _T_274 ? _GEN_3 : _T_718_17;
  assign _GEN_247 = 5'h12 == _T_274 ? _GEN_3 : _T_718_18;
  assign _GEN_248 = 5'h13 == _T_274 ? _GEN_3 : _T_718_19;
  assign _GEN_249 = 5'h14 == _T_274 ? _GEN_3 : _T_718_20;
  assign _GEN_250 = 5'h15 == _T_274 ? _GEN_3 : _T_718_21;
  assign _GEN_251 = 5'h16 == _T_274 ? _GEN_3 : _T_718_22;
  assign _GEN_252 = 5'h17 == _T_274 ? _GEN_3 : _T_718_23;
  assign _GEN_253 = 5'h18 == _T_274 ? _GEN_3 : _T_718_24;
  assign _GEN_254 = 5'h19 == _T_274 ? _GEN_3 : _T_718_25;
  assign _GEN_255 = 5'h1a == _T_274 ? _GEN_3 : _T_718_26;
  assign _GEN_256 = 5'h1b == _T_274 ? _GEN_3 : _T_718_27;
  assign _GEN_257 = 5'h1c == _T_274 ? _GEN_3 : _T_718_28;
  assign _GEN_258 = 5'h1d == _T_274 ? _GEN_3 : _T_718_29;
  assign _GEN_259 = 5'h1e == _T_274 ? _GEN_3 : _T_718_30;
  assign _GEN_260 = 5'h1f == _T_274 ? _GEN_3 : _T_718_31;
  assign _GEN_261 = _T_764 ? _GEN_229 : _T_718_0;
  assign _GEN_262 = _T_764 ? _GEN_230 : _T_718_1;
  assign _GEN_263 = _T_764 ? _GEN_231 : _T_718_2;
  assign _GEN_264 = _T_764 ? _GEN_232 : _T_718_3;
  assign _GEN_265 = _T_764 ? _GEN_233 : _T_718_4;
  assign _GEN_266 = _T_764 ? _GEN_234 : _T_718_5;
  assign _GEN_267 = _T_764 ? _GEN_235 : _T_718_6;
  assign _GEN_268 = _T_764 ? _GEN_236 : _T_718_7;
  assign _GEN_269 = _T_764 ? _GEN_237 : _T_718_8;
  assign _GEN_270 = _T_764 ? _GEN_238 : _T_718_9;
  assign _GEN_271 = _T_764 ? _GEN_239 : _T_718_10;
  assign _GEN_272 = _T_764 ? _GEN_240 : _T_718_11;
  assign _GEN_273 = _T_764 ? _GEN_241 : _T_718_12;
  assign _GEN_274 = _T_764 ? _GEN_242 : _T_718_13;
  assign _GEN_275 = _T_764 ? _GEN_243 : _T_718_14;
  assign _GEN_276 = _T_764 ? _GEN_244 : _T_718_15;
  assign _GEN_277 = _T_764 ? _GEN_245 : _T_718_16;
  assign _GEN_278 = _T_764 ? _GEN_246 : _T_718_17;
  assign _GEN_279 = _T_764 ? _GEN_247 : _T_718_18;
  assign _GEN_280 = _T_764 ? _GEN_248 : _T_718_19;
  assign _GEN_281 = _T_764 ? _GEN_249 : _T_718_20;
  assign _GEN_282 = _T_764 ? _GEN_250 : _T_718_21;
  assign _GEN_283 = _T_764 ? _GEN_251 : _T_718_22;
  assign _GEN_284 = _T_764 ? _GEN_252 : _T_718_23;
  assign _GEN_285 = _T_764 ? _GEN_253 : _T_718_24;
  assign _GEN_286 = _T_764 ? _GEN_254 : _T_718_25;
  assign _GEN_287 = _T_764 ? _GEN_255 : _T_718_26;
  assign _GEN_288 = _T_764 ? _GEN_256 : _T_718_27;
  assign _GEN_289 = _T_764 ? _GEN_257 : _T_718_28;
  assign _GEN_290 = _T_764 ? _GEN_258 : _T_718_29;
  assign _GEN_291 = _T_764 ? _GEN_259 : _T_718_30;
  assign _GEN_292 = _T_764 ? _GEN_260 : _T_718_31;
  assign _T_768 = _T_703 & _T_268;
  assign _T_770 = _T_714 == 1'h0;
  assign _T_771 = _T_768 & _T_770;
  assign _GEN_293 = _T_771 ? 1'h1 : _T_711;
  assign _T_773 = _T_711 & io_outputMemAddrReadys_1;
  assign _GEN_294 = _T_773 ? 1'h0 : _GEN_293;
  assign _GEN_295 = _T_773 ? 1'h1 : _T_714;
  assign _T_776 = {_T_718_1,_T_718_0};
  assign _T_777 = {_T_718_3,_T_718_2};
  assign _T_778 = {_T_777,_T_776};
  assign _T_779 = {_T_718_5,_T_718_4};
  assign _T_780 = {_T_718_7,_T_718_6};
  assign _T_781 = {_T_780,_T_779};
  assign _T_782 = {_T_781,_T_778};
  assign _T_783 = {_T_718_9,_T_718_8};
  assign _T_784 = {_T_718_11,_T_718_10};
  assign _T_785 = {_T_784,_T_783};
  assign _T_786 = {_T_718_13,_T_718_12};
  assign _T_787 = {_T_718_15,_T_718_14};
  assign _T_788 = {_T_787,_T_786};
  assign _T_789 = {_T_788,_T_785};
  assign _T_790 = {_T_789,_T_782};
  assign _T_791 = {_T_718_17,_T_718_16};
  assign _T_792 = {_T_718_19,_T_718_18};
  assign _T_793 = {_T_792,_T_791};
  assign _T_794 = {_T_718_21,_T_718_20};
  assign _T_795 = {_T_718_23,_T_718_22};
  assign _T_796 = {_T_795,_T_794};
  assign _T_797 = {_T_796,_T_793};
  assign _T_798 = {_T_718_25,_T_718_24};
  assign _T_799 = {_T_718_27,_T_718_26};
  assign _T_800 = {_T_799,_T_798};
  assign _T_801 = {_T_718_29,_T_718_28};
  assign _T_802 = {_T_718_31,_T_718_30};
  assign _T_803 = {_T_802,_T_801};
  assign _T_804 = {_T_803,_T_800};
  assign _T_805 = {_T_804,_T_797};
  assign _T_806 = {_T_805,_T_790};
  assign _T_810 = _T_288 ? io_outputMemAddrReadys_1 : 1'h0;
  assign _T_813 = io_outputMemBlockReadys_1 & _T_755;
  assign _T_815 = _T_288 ? _T_813 : 1'h0;
  assign _T_816 = io_outputMemBlockReadys_1 & io_outputMemBlockValids_1;
  assign _T_823 = _T_276 | _T_813;
  assign _T_824 = _T_703 & _T_823;
  assign _T_829 = _T_288 + 1'h1;
  assign _T_830 = _T_829[0:0];
  assign _T_831 = _T_288 ? 1'h1 : _T_830;
  assign _GEN_296 = _T_824 ? _T_831 : _T_288;
  assign _GEN_297 = _T_824 ? 1'h0 : _GEN_228;
  assign _GEN_298 = _T_824 ? 1'h0 : _GEN_227;
  assign _GEN_299 = _T_824 ? 1'h0 : _GEN_295;
  assign cumFinished = cores_0_outputFinished & cores_1_outputFinished;
  assign io_inputMemAddrs_0 = _T_238;
  assign io_inputMemAddrs_1 = _T_246;
  assign io_inputMemAddrValids_0 = _T_299;
  assign io_inputMemAddrValids_1 = _T_438;
  assign io_inputMemBlockReadys_0 = _T_403;
  assign io_inputMemBlockReadys_1 = _T_542;
  assign io_outputMemAddrs_0 = _T_254;
  assign io_outputMemAddrs_1 = _T_266;
  assign io_outputMemAddrValids_0 = _T_577;
  assign io_outputMemAddrValids_1 = _T_711;
  assign io_outputMemBlocks_0 = _T_672;
  assign io_outputMemBlocks_1 = _T_806;
  assign io_outputMemBlockValids_0 = _T_621;
  assign io_outputMemBlockValids_1 = _T_755;
  assign io_finished = cumFinished;
  assign StreamingCore_io_inputMemAddrReady = cores_0_inputMemAddrReady;
  assign StreamingCore_io_inputMemBlock = cores_0_inputMemBlock;
  assign StreamingCore_io_inputMemIdx = cores_0_inputMemIdx;
  assign StreamingCore_io_inputMemBlockValid = cores_0_inputMemBlockValid;
  assign StreamingCore_io_outputMemAddrReady = cores_0_outputMemAddrReady;
  assign StreamingCore_io_outputMemBlockReady = cores_0_outputMemBlockReady;
  assign StreamingCore_clock = clock;
  assign StreamingCore_reset = reset;
  assign StreamingCore_1_io_inputMemAddrReady = cores_1_inputMemAddrReady;
  assign StreamingCore_1_io_inputMemBlock = cores_1_inputMemBlock;
  assign StreamingCore_1_io_inputMemIdx = cores_1_inputMemIdx;
  assign StreamingCore_1_io_inputMemBlockValid = cores_1_inputMemBlockValid;
  assign StreamingCore_1_io_outputMemAddrReady = cores_1_outputMemAddrReady;
  assign StreamingCore_1_io_outputMemBlockReady = cores_1_outputMemBlockReady;
  assign StreamingCore_1_clock = clock;
  assign StreamingCore_1_reset = reset;
  assign cores_0_inputMemAddr = StreamingCore_io_inputMemAddr;
  assign cores_0_inputMemAddrValid = StreamingCore_io_inputMemAddrValid;
  assign cores_0_inputMemAddrReady = _T_407;
  assign cores_0_inputMemBlock = _GEN_0;
  assign cores_0_inputMemIdx = _T_343;
  assign cores_0_inputMemBlockValid = _T_412;
  assign cores_0_inputMemBlockReady = StreamingCore_io_inputMemBlockReady;
  assign cores_0_outputMemAddr = StreamingCore_io_outputMemAddr;
  assign cores_0_outputMemAddrValid = StreamingCore_io_outputMemAddrValid;
  assign cores_0_outputMemAddrReady = _T_676;
  assign cores_0_outputMemBlock = StreamingCore_io_outputMemBlock;
  assign cores_0_outputMemIdx = StreamingCore_io_outputMemIdx;
  assign cores_0_outputMemBlockValid = StreamingCore_io_outputMemBlockValid;
  assign cores_0_outputMemBlockReady = _T_681;
  assign cores_0_inputFinished = StreamingCore_io_inputFinished;
  assign cores_0_outputFinished = StreamingCore_io_outputFinished;
  assign cores_1_inputMemAddr = StreamingCore_1_io_inputMemAddr;
  assign cores_1_inputMemAddrValid = StreamingCore_1_io_inputMemAddrValid;
  assign cores_1_inputMemAddrReady = _T_546;
  assign cores_1_inputMemBlock = _GEN_1;
  assign cores_1_inputMemIdx = _T_482;
  assign cores_1_inputMemBlockValid = _T_551;
  assign cores_1_inputMemBlockReady = StreamingCore_1_io_inputMemBlockReady;
  assign cores_1_outputMemAddr = StreamingCore_1_io_outputMemAddr;
  assign cores_1_outputMemAddrValid = StreamingCore_1_io_outputMemAddrValid;
  assign cores_1_outputMemAddrReady = _T_810;
  assign cores_1_outputMemBlock = StreamingCore_1_io_outputMemBlock;
  assign cores_1_outputMemIdx = StreamingCore_1_io_outputMemIdx;
  assign cores_1_outputMemBlockValid = StreamingCore_1_io_outputMemBlockValid;
  assign cores_1_outputMemBlockReady = _T_815;
  assign cores_1_inputFinished = StreamingCore_1_io_inputFinished;
  assign cores_1_outputFinished = StreamingCore_1_io_outputFinished;
  assign _GEN_0 = _GEN_75;
  assign _GEN_1 = _GEN_150;
  assign _GEN_2 = _T_260;
  assign _GEN_3 = _T_272;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{$random}};
  _T_238 = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_240 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_242 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_244 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{$random}};
  _T_246 = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_248 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_250 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_252 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{$random}};
  _T_254 = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_256 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_258 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_260 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_262 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_264 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{$random}};
  _T_266 = _RAND_14[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_268 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_270 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_272 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_274 = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_276 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_279 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_282 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_285 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_288 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_291 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_299 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_302 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_306_0 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_306_1 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_306_2 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_306_3 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_306_4 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_306_5 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_306_6 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_306_7 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_306_8 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_306_9 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_306_10 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_306_11 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_306_12 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_306_13 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_306_14 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_306_15 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_306_16 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_306_17 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_306_18 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_306_19 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_306_20 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_306_21 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_306_22 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_306_23 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_306_24 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_306_25 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_306_26 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_306_27 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_306_28 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_306_29 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_306_30 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_306_31 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_343 = _RAND_59[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_346 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_430 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_438 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_441 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_445_0 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_445_1 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_445_2 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_445_3 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_445_4 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_445_5 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_445_6 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_445_7 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_445_8 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_445_9 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_445_10 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_445_11 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_445_12 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_445_13 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_445_14 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_445_15 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_445_16 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_445_17 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_445_18 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_445_19 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_445_20 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_445_21 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_445_22 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_445_23 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_445_24 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_445_25 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_445_26 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_445_27 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_445_28 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_445_29 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_445_30 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_445_31 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_482 = _RAND_96[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_485 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_569 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_577 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_580 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_584_0 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_584_1 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_584_2 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_584_3 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_584_4 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_584_5 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_584_6 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_584_7 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_584_8 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_584_9 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_584_10 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_584_11 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_584_12 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_584_13 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_584_14 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_584_15 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_584_16 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_584_17 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_584_18 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_584_19 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_584_20 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_584_21 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_584_22 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_584_23 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_584_24 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_584_25 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_584_26 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_584_27 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_584_28 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_584_29 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_584_30 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_584_31 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_621 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_703 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  _T_711 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_714 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  _T_718_0 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  _T_718_1 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  _T_718_2 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  _T_718_3 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  _T_718_4 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  _T_718_5 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  _T_718_6 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  _T_718_7 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  _T_718_8 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  _T_718_9 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  _T_718_10 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  _T_718_11 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  _T_718_12 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  _T_718_13 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  _T_718_14 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  _T_718_15 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  _T_718_16 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  _T_718_17 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _T_718_18 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  _T_718_19 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _T_718_20 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  _T_718_21 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  _T_718_22 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _T_718_23 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  _T_718_24 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  _T_718_25 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  _T_718_26 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  _T_718_27 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  _T_718_28 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  _T_718_29 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  _T_718_30 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  _T_718_31 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  _T_755 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_238 <= cores_0_inputMemAddr;
    _T_240 <= cores_0_inputMemAddrValid;
    _T_242 <= cores_0_inputMemBlockReady;
    _T_244 <= cores_0_inputFinished;
    _T_246 <= cores_1_inputMemAddr;
    _T_248 <= cores_1_inputMemAddrValid;
    _T_250 <= cores_1_inputMemBlockReady;
    _T_252 <= cores_1_inputFinished;
    _T_254 <= cores_0_outputMemAddr;
    _T_256 <= cores_0_outputMemAddrValid;
    _T_258 <= cores_0_outputMemBlockValid;
    _T_260 <= cores_0_outputMemBlock;
    _T_262 <= cores_0_outputMemIdx;
    _T_264 <= cores_0_outputFinished;
    _T_266 <= cores_1_outputMemAddr;
    _T_268 <= cores_1_outputMemAddrValid;
    _T_270 <= cores_1_outputMemBlockValid;
    _T_272 <= cores_1_outputMemBlock;
    _T_274 <= cores_1_outputMemIdx;
    _T_276 <= cores_1_outputFinished;
    if (reset) begin
      _T_279 <= 1'h0;
    end else begin
      if (_T_418) begin
        if (_T_405) begin
          _T_279 <= 1'h0;
        end else begin
          _T_279 <= _T_424;
        end
      end
    end
    if (reset) begin
      _T_282 <= 1'h1;
    end else begin
      if (_T_557) begin
        if (_T_282) begin
          _T_282 <= 1'h1;
        end else begin
          _T_282 <= _T_563;
        end
      end
    end
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (_T_674) begin
          _T_285 <= 1'h0;
        end else begin
          _T_285 <= _T_696;
        end
      end
    end
    if (reset) begin
      _T_288 <= 1'h1;
    end else begin
      if (_T_824) begin
        if (_T_288) begin
          _T_288 <= 1'h1;
        end else begin
          _T_288 <= _T_830;
        end
      end
    end
    if (reset) begin
      _T_291 <= 1'h0;
    end else begin
      if (_T_418) begin
        _T_291 <= 1'h0;
      end else begin
        if (_T_293) begin
          _T_291 <= _T_296;
        end
      end
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      if (_T_398) begin
        _T_299 <= 1'h0;
      end else begin
        if (_T_396) begin
          _T_299 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_302 <= 1'h0;
    end else begin
      if (_T_418) begin
        _T_302 <= 1'h0;
      end else begin
        if (_T_398) begin
          _T_302 <= 1'h1;
        end
      end
    end
    if (_T_347) begin
      _T_306_0 <= _T_348;
    end
    if (_T_347) begin
      _T_306_1 <= _T_349;
    end
    if (_T_347) begin
      _T_306_2 <= _T_350;
    end
    if (_T_347) begin
      _T_306_3 <= _T_351;
    end
    if (_T_347) begin
      _T_306_4 <= _T_352;
    end
    if (_T_347) begin
      _T_306_5 <= _T_353;
    end
    if (_T_347) begin
      _T_306_6 <= _T_354;
    end
    if (_T_347) begin
      _T_306_7 <= _T_355;
    end
    if (_T_347) begin
      _T_306_8 <= _T_356;
    end
    if (_T_347) begin
      _T_306_9 <= _T_357;
    end
    if (_T_347) begin
      _T_306_10 <= _T_358;
    end
    if (_T_347) begin
      _T_306_11 <= _T_359;
    end
    if (_T_347) begin
      _T_306_12 <= _T_360;
    end
    if (_T_347) begin
      _T_306_13 <= _T_361;
    end
    if (_T_347) begin
      _T_306_14 <= _T_362;
    end
    if (_T_347) begin
      _T_306_15 <= _T_363;
    end
    if (_T_347) begin
      _T_306_16 <= _T_364;
    end
    if (_T_347) begin
      _T_306_17 <= _T_365;
    end
    if (_T_347) begin
      _T_306_18 <= _T_366;
    end
    if (_T_347) begin
      _T_306_19 <= _T_367;
    end
    if (_T_347) begin
      _T_306_20 <= _T_368;
    end
    if (_T_347) begin
      _T_306_21 <= _T_369;
    end
    if (_T_347) begin
      _T_306_22 <= _T_370;
    end
    if (_T_347) begin
      _T_306_23 <= _T_371;
    end
    if (_T_347) begin
      _T_306_24 <= _T_372;
    end
    if (_T_347) begin
      _T_306_25 <= _T_373;
    end
    if (_T_347) begin
      _T_306_26 <= _T_374;
    end
    if (_T_347) begin
      _T_306_27 <= _T_375;
    end
    if (_T_347) begin
      _T_306_28 <= _T_376;
    end
    if (_T_347) begin
      _T_306_29 <= _T_377;
    end
    if (_T_347) begin
      _T_306_30 <= _T_378;
    end
    if (_T_347) begin
      _T_306_31 <= _T_379;
    end
    if (reset) begin
      _T_343 <= 5'h0;
    end else begin
      if (_T_346) begin
        if (_T_385) begin
          _T_343 <= 5'h0;
        end else begin
          _T_343 <= _T_390;
        end
      end
    end
    if (reset) begin
      _T_346 <= 1'h0;
    end else begin
      if (_T_346) begin
        if (_T_385) begin
          _T_346 <= 1'h0;
        end else begin
          if (_T_347) begin
            _T_346 <= 1'h1;
          end
        end
      end else begin
        if (_T_347) begin
          _T_346 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_430 <= 1'h0;
    end else begin
      if (_T_557) begin
        _T_430 <= 1'h0;
      end else begin
        if (_T_432) begin
          _T_430 <= _T_435;
        end
      end
    end
    if (reset) begin
      _T_438 <= 1'h0;
    end else begin
      if (_T_537) begin
        _T_438 <= 1'h0;
      end else begin
        if (_T_535) begin
          _T_438 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_441 <= 1'h0;
    end else begin
      if (_T_557) begin
        _T_441 <= 1'h0;
      end else begin
        if (_T_537) begin
          _T_441 <= 1'h1;
        end
      end
    end
    if (_T_486) begin
      _T_445_0 <= _T_487;
    end
    if (_T_486) begin
      _T_445_1 <= _T_488;
    end
    if (_T_486) begin
      _T_445_2 <= _T_489;
    end
    if (_T_486) begin
      _T_445_3 <= _T_490;
    end
    if (_T_486) begin
      _T_445_4 <= _T_491;
    end
    if (_T_486) begin
      _T_445_5 <= _T_492;
    end
    if (_T_486) begin
      _T_445_6 <= _T_493;
    end
    if (_T_486) begin
      _T_445_7 <= _T_494;
    end
    if (_T_486) begin
      _T_445_8 <= _T_495;
    end
    if (_T_486) begin
      _T_445_9 <= _T_496;
    end
    if (_T_486) begin
      _T_445_10 <= _T_497;
    end
    if (_T_486) begin
      _T_445_11 <= _T_498;
    end
    if (_T_486) begin
      _T_445_12 <= _T_499;
    end
    if (_T_486) begin
      _T_445_13 <= _T_500;
    end
    if (_T_486) begin
      _T_445_14 <= _T_501;
    end
    if (_T_486) begin
      _T_445_15 <= _T_502;
    end
    if (_T_486) begin
      _T_445_16 <= _T_503;
    end
    if (_T_486) begin
      _T_445_17 <= _T_504;
    end
    if (_T_486) begin
      _T_445_18 <= _T_505;
    end
    if (_T_486) begin
      _T_445_19 <= _T_506;
    end
    if (_T_486) begin
      _T_445_20 <= _T_507;
    end
    if (_T_486) begin
      _T_445_21 <= _T_508;
    end
    if (_T_486) begin
      _T_445_22 <= _T_509;
    end
    if (_T_486) begin
      _T_445_23 <= _T_510;
    end
    if (_T_486) begin
      _T_445_24 <= _T_511;
    end
    if (_T_486) begin
      _T_445_25 <= _T_512;
    end
    if (_T_486) begin
      _T_445_26 <= _T_513;
    end
    if (_T_486) begin
      _T_445_27 <= _T_514;
    end
    if (_T_486) begin
      _T_445_28 <= _T_515;
    end
    if (_T_486) begin
      _T_445_29 <= _T_516;
    end
    if (_T_486) begin
      _T_445_30 <= _T_517;
    end
    if (_T_486) begin
      _T_445_31 <= _T_518;
    end
    if (reset) begin
      _T_482 <= 5'h0;
    end else begin
      if (_T_485) begin
        if (_T_524) begin
          _T_482 <= 5'h0;
        end else begin
          _T_482 <= _T_529;
        end
      end
    end
    if (reset) begin
      _T_485 <= 1'h0;
    end else begin
      if (_T_485) begin
        if (_T_524) begin
          _T_485 <= 1'h0;
        end else begin
          if (_T_486) begin
            _T_485 <= 1'h1;
          end
        end
      end else begin
        if (_T_486) begin
          _T_485 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_569 <= 1'h0;
    end else begin
      if (_T_690) begin
        _T_569 <= 1'h0;
      end else begin
        if (_T_571) begin
          _T_569 <= _T_574;
        end
      end
    end
    if (reset) begin
      _T_577 <= 1'h0;
    end else begin
      if (_T_639) begin
        _T_577 <= 1'h0;
      end else begin
        if (_T_637) begin
          _T_577 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_580 <= 1'h0;
    end else begin
      if (_T_690) begin
        _T_580 <= 1'h0;
      end else begin
        if (_T_639) begin
          _T_580 <= 1'h1;
        end
      end
    end
    if (_T_630) begin
      if (5'h0 == _T_262) begin
        _T_584_0 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h1 == _T_262) begin
        _T_584_1 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h2 == _T_262) begin
        _T_584_2 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h3 == _T_262) begin
        _T_584_3 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h4 == _T_262) begin
        _T_584_4 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h5 == _T_262) begin
        _T_584_5 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h6 == _T_262) begin
        _T_584_6 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h7 == _T_262) begin
        _T_584_7 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h8 == _T_262) begin
        _T_584_8 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h9 == _T_262) begin
        _T_584_9 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'ha == _T_262) begin
        _T_584_10 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'hb == _T_262) begin
        _T_584_11 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'hc == _T_262) begin
        _T_584_12 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'hd == _T_262) begin
        _T_584_13 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'he == _T_262) begin
        _T_584_14 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'hf == _T_262) begin
        _T_584_15 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h10 == _T_262) begin
        _T_584_16 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h11 == _T_262) begin
        _T_584_17 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h12 == _T_262) begin
        _T_584_18 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h13 == _T_262) begin
        _T_584_19 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h14 == _T_262) begin
        _T_584_20 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h15 == _T_262) begin
        _T_584_21 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h16 == _T_262) begin
        _T_584_22 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h17 == _T_262) begin
        _T_584_23 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h18 == _T_262) begin
        _T_584_24 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h19 == _T_262) begin
        _T_584_25 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h1a == _T_262) begin
        _T_584_26 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h1b == _T_262) begin
        _T_584_27 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h1c == _T_262) begin
        _T_584_28 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h1d == _T_262) begin
        _T_584_29 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h1e == _T_262) begin
        _T_584_30 <= _GEN_2;
      end
    end
    if (_T_630) begin
      if (5'h1f == _T_262) begin
        _T_584_31 <= _GEN_2;
      end
    end
    if (reset) begin
      _T_621 <= 1'h0;
    end else begin
      if (_T_690) begin
        _T_621 <= 1'h0;
      end else begin
        if (_T_627) begin
          _T_621 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_703 <= 1'h0;
    end else begin
      if (_T_824) begin
        _T_703 <= 1'h0;
      end else begin
        if (_T_705) begin
          _T_703 <= _T_708;
        end
      end
    end
    if (reset) begin
      _T_711 <= 1'h0;
    end else begin
      if (_T_773) begin
        _T_711 <= 1'h0;
      end else begin
        if (_T_771) begin
          _T_711 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_714 <= 1'h0;
    end else begin
      if (_T_824) begin
        _T_714 <= 1'h0;
      end else begin
        if (_T_773) begin
          _T_714 <= 1'h1;
        end
      end
    end
    if (_T_764) begin
      if (5'h0 == _T_274) begin
        _T_718_0 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h1 == _T_274) begin
        _T_718_1 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h2 == _T_274) begin
        _T_718_2 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h3 == _T_274) begin
        _T_718_3 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h4 == _T_274) begin
        _T_718_4 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h5 == _T_274) begin
        _T_718_5 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h6 == _T_274) begin
        _T_718_6 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h7 == _T_274) begin
        _T_718_7 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h8 == _T_274) begin
        _T_718_8 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h9 == _T_274) begin
        _T_718_9 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'ha == _T_274) begin
        _T_718_10 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'hb == _T_274) begin
        _T_718_11 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'hc == _T_274) begin
        _T_718_12 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'hd == _T_274) begin
        _T_718_13 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'he == _T_274) begin
        _T_718_14 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'hf == _T_274) begin
        _T_718_15 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h10 == _T_274) begin
        _T_718_16 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h11 == _T_274) begin
        _T_718_17 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h12 == _T_274) begin
        _T_718_18 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h13 == _T_274) begin
        _T_718_19 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h14 == _T_274) begin
        _T_718_20 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h15 == _T_274) begin
        _T_718_21 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h16 == _T_274) begin
        _T_718_22 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h17 == _T_274) begin
        _T_718_23 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h18 == _T_274) begin
        _T_718_24 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h19 == _T_274) begin
        _T_718_25 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h1a == _T_274) begin
        _T_718_26 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h1b == _T_274) begin
        _T_718_27 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h1c == _T_274) begin
        _T_718_28 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h1d == _T_274) begin
        _T_718_29 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h1e == _T_274) begin
        _T_718_30 <= _GEN_3;
      end
    end
    if (_T_764) begin
      if (5'h1f == _T_274) begin
        _T_718_31 <= _GEN_3;
      end
    end
    if (reset) begin
      _T_755 <= 1'h0;
    end else begin
      if (_T_824) begin
        _T_755 <= 1'h0;
      end else begin
        if (_T_761) begin
          _T_755 <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_347 & _T_383) begin
          $fwrite(32'h80000002,"inputBuffer: 0x%h for core %d, channel 0\n",io_inputMemBlocks_0,_T_279);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_486 & _T_383) begin
          $fwrite(32'h80000002,"inputBuffer: 0x%h for core %d, channel 1\n",io_inputMemBlocks_1,_T_282);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_682 & _T_383) begin
          $fwrite(32'h80000002,"outputBuffer: 0x%h for core %d, channel 0\n",io_outputMemBlocks_0,_T_285);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_816 & _T_383) begin
          $fwrite(32'h80000002,"outputBuffer: 0x%h for core %d, channel 1\n",io_outputMemBlocks_1,_T_288);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
