// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

module cl_hello_world 

(
   `include "cl_ports.vh" // Fixed port definition

);

`include "cl_common_defines.vh"      // CL Defines for all examples
`include "cl_id_defines.vh"          // Defines for ID0 and ID1 (PCI ID's)
`include "cl_hello_world_defines.vh" // CL Defines for cl_hello_world

logic rst_main_n_sync;


//--------------------------------------------0
// Start with Tie-Off of Unused Interfaces
//---------------------------------------------
// the developer should use the next set of `include
// to properly tie-off any unused interface
// The list is put in the top of the module
// to avoid cases where developer may forget to
// remove it from the end of the file

// `include "unused_flr_template.inc"
`include "unused_ddr_a_b_d_template.inc"
`include "unused_ddr_c_template.inc"
`include "unused_pcim_template.inc"
// `include "unused_dma_pcis_template.inc"
`include "unused_cl_sda_template.inc"
`include "unused_sh_bar1_template.inc"
`include "unused_apppf_irq_template.inc"
`include "unused_hmc_template.inc"
`include "unused_aurora_template.inc"

//-------------------------------------------------
// Wires
//-------------------------------------------------
  logic        arvalid_q;
  logic [31:0] araddr_q;
  logic [31:0] hello_world_q_byte_swapped;
  logic [15:0] vled_q;
  logic [15:0] pre_cl_sh_status_vled;
  logic [15:0] sh_cl_status_vdip_q;
  logic [15:0] sh_cl_status_vdip_q2;
  logic [31:0] hello_world_q;

//-------------------------------------------------
// ID Values (cl_hello_world_defines.vh)
//-------------------------------------------------
  assign cl_sh_id0[31:0] = `CL_SH_ID0;
  assign cl_sh_id1[31:0] = `CL_SH_ID1;

//-------------------------------------------------
// Reset Synchronization
//-------------------------------------------------
logic pre_sync_rst_n;

always_ff @(negedge rst_main_n or posedge clk_main_a0)
   if (!rst_main_n)
   begin
      pre_sync_rst_n  <= 0;
      rst_main_n_sync <= 0;
   end
   else
   begin
      pre_sync_rst_n  <= 1;
      rst_main_n_sync <= pre_sync_rst_n;
   end

//-------------------------------------------------
// PCIe OCL AXI-L (SH to CL) Timing Flops
//-------------------------------------------------

  // Write address                                                                                                              
  logic        sh_ocl_awvalid_q;
  logic [31:0] sh_ocl_awaddr_q;
  logic        ocl_sh_awready_q;
                                                                                                                              
  // Write data                                                                                                                
  logic        sh_ocl_wvalid_q;
  logic [31:0] sh_ocl_wdata_q;
  logic [ 3:0] sh_ocl_wstrb_q;
  logic        ocl_sh_wready_q;
                                                                                                                              
  // Write response                                                                                                            
  logic        ocl_sh_bvalid_q;
  logic [ 1:0] ocl_sh_bresp_q;
  logic        sh_ocl_bready_q;
                                                                                                                              
  // Read address                                                                                                              
  logic        sh_ocl_arvalid_q;
  logic [31:0] sh_ocl_araddr_q;
  logic        ocl_sh_arready_q;
                                                                                                                              
  // Read data/response                                                                                                        
  logic        ocl_sh_rvalid_q;
  logic [31:0] ocl_sh_rdata_q;
  logic [ 1:0] ocl_sh_rresp_q;
  logic        sh_ocl_rready_q;

/*
  axi_register_slice_light AXIL_OCL_REG_SLC (
   .aclk          (clk_main_a0),
   .aresetn       (rst_main_n_sync),
   .s_axi_awaddr  (sh_ocl_awaddr),
   .s_axi_awprot   (2'h0),
   .s_axi_awvalid (sh_ocl_awvalid),
   .s_axi_awready (ocl_sh_awready),
   .s_axi_wdata   (sh_ocl_wdata),
   .s_axi_wstrb   (sh_ocl_wstrb),
   .s_axi_wvalid  (sh_ocl_wvalid),
   .s_axi_wready  (ocl_sh_wready),
   .s_axi_bresp   (ocl_sh_bresp),
   .s_axi_bvalid  (ocl_sh_bvalid),
   .s_axi_bready  (sh_ocl_bready),
   .s_axi_araddr  (sh_ocl_araddr),
   .s_axi_arvalid (sh_ocl_arvalid),
   .s_axi_arready (ocl_sh_arready),
   .s_axi_rdata   (ocl_sh_rdata),
   .s_axi_rresp   (ocl_sh_rresp),
   .s_axi_rvalid  (ocl_sh_rvalid),
   .s_axi_rready  (sh_ocl_rready),
   .m_axi_awaddr  (sh_ocl_awaddr_q),
   .m_axi_awprot  (),
   .m_axi_awvalid (sh_ocl_awvalid_q),
   .m_axi_awready (ocl_sh_awready_q),
   .m_axi_wdata   (sh_ocl_wdata_q),
   .m_axi_wstrb   (sh_ocl_wstrb_q),
   .m_axi_wvalid  (sh_ocl_wvalid_q),
   .m_axi_wready  (ocl_sh_wready_q),
   .m_axi_bresp   (ocl_sh_bresp_q),
   .m_axi_bvalid  (ocl_sh_bvalid_q),
   .m_axi_bready  (sh_ocl_bready_q),
   .m_axi_araddr  (sh_ocl_araddr_q),
   .m_axi_arvalid (sh_ocl_arvalid_q),
   .m_axi_arready (ocl_sh_arready_q),
   .m_axi_rdata   (ocl_sh_rdata_q),
   .m_axi_rresp   (ocl_sh_rresp_q),
   .m_axi_rvalid  (ocl_sh_rvalid_q),
   .m_axi_rready  (sh_ocl_rready_q)
  );

//--------------------------------------------------------------
// PCIe OCL AXI-L Slave Accesses (accesses from PCIe AppPF BAR0)
//--------------------------------------------------------------
// Only supports single-beat accesses.

   logic        awvalid;
   logic [31:0] awaddr;
   logic        wvalid;
   logic [31:0] wdata;
   logic [3:0]  wstrb;
   logic        bready;
   logic        arvalid;
   logic [31:0] araddr;
   logic        rready;

   logic        awready;
   logic        wready;
   logic        bvalid;
   logic [1:0]  bresp;
   logic        arready;
   logic        rvalid;
   logic [31:0] rdata;
   logic [1:0]  rresp;

   // Inputs
   assign awvalid         = sh_ocl_awvalid_q;
   assign awaddr[31:0]    = sh_ocl_awaddr_q;
   assign wvalid          = sh_ocl_wvalid_q;
   assign wdata[31:0]     = sh_ocl_wdata_q;
   assign wstrb[3:0]      = sh_ocl_wstrb_q;
   assign bready          = sh_ocl_bready_q;
   assign arvalid         = sh_ocl_arvalid_q;
   assign araddr[31:0]    = sh_ocl_araddr_q;
   assign rready          = sh_ocl_rready_q;

   // Outputs
   assign ocl_sh_awready_q = awready;
   assign ocl_sh_wready_q  = wready;
   assign ocl_sh_bvalid_q  = bvalid;
   assign ocl_sh_bresp_q   = bresp[1:0];
   assign ocl_sh_arready_q = arready;
   assign ocl_sh_rvalid_q  = rvalid;
   assign ocl_sh_rdata_q   = rdata;
   assign ocl_sh_rresp_q   = rresp[1:0];

// Write Request
logic        wr_active;
logic [31:0] wr_addr;

always_ff @(posedge clk_main_a0)
  if (!rst_main_n_sync) begin
     wr_active <= 0;
     wr_addr   <= 0;
  end
  else begin
     wr_active <=  wr_active && bvalid  && bready ? 1'b0     :
                  ~wr_active && awvalid           ? 1'b1     :
                                                    wr_active;
     wr_addr <= awvalid && ~wr_active ? awaddr : wr_addr     ;
  end

assign awready = ~wr_active;
assign wready  =  wr_active && wvalid;

// Write Response
always_ff @(posedge clk_main_a0)
  if (!rst_main_n_sync) 
    bvalid <= 0;
  else
    bvalid <=  bvalid &&  bready           ? 1'b0  : 
                         ~bvalid && wready ? 1'b1  :
                                             bvalid;
assign bresp = 0;

// Read Request
always_ff @(posedge clk_main_a0)
   if (!rst_main_n_sync) begin
      arvalid_q <= 0;
      araddr_q  <= 0;
   end
   else begin
      arvalid_q <= arvalid;
      araddr_q  <= arvalid ? araddr : araddr_q;
   end

assign arready = !arvalid_q && !rvalid;

// Read Response
always_ff @(posedge clk_main_a0)
   if (!rst_main_n_sync)
   begin
      rvalid <= 0;
      rdata  <= 0;
      rresp  <= 0;
   end
   else if (rvalid && rready)
   begin
      rvalid <= 0;
      rdata  <= 0;
      rresp  <= 0;
   end
   else if (arvalid_q) 
   begin
      rvalid <= 1;
      rdata  <= (araddr_q == `HELLO_WORLD_REG_ADDR) ? hello_world_q_byte_swapped[31:0]:
                (araddr_q == `VLED_REG_ADDR       ) ? {16'b0,vled_q[15:0]            }:
                                                      `UNIMPLEMENTED_REG_VALUE        ;
      rresp  <= 0;
   end
*/

axi_register_slice PCI_AXL_REG_SLC (
    .aclk          (clk_main_a0),
    .aresetn       (!rst_main_n_sync),
    .s_axi_awid    (sh_cl_dma_pcis_bus.awid),
    .s_axi_awaddr  (sh_cl_dma_pcis_bus.awaddr),
    .s_axi_awlen   (sh_cl_dma_pcis_bus.awlen),                                            
    .s_axi_awvalid (sh_cl_dma_pcis_bus.awvalid),
    .s_axi_awsize  (sh_cl_dma_pcis_bus.awsize),
    .s_axi_awready (sh_cl_dma_pcis_bus.awready),
    .s_axi_wdata   (sh_cl_dma_pcis_bus.wdata),
    .s_axi_wstrb   (sh_cl_dma_pcis_bus.wstrb),
    .s_axi_wlast   (sh_cl_dma_pcis_bus.wlast),
    .s_axi_wvalid  (sh_cl_dma_pcis_bus.wvalid),
    .s_axi_wready  (sh_cl_dma_pcis_bus.wready),
    .s_axi_bid     (sh_cl_dma_pcis_bus.bid),
    .s_axi_bresp   (sh_cl_dma_pcis_bus.bresp),
    .s_axi_bvalid  (sh_cl_dma_pcis_bus.bvalid),
    .s_axi_bready  (sh_cl_dma_pcis_bus.bready),
    .s_axi_arid    (sh_cl_dma_pcis_bus.arid),
    .s_axi_araddr  (sh_cl_dma_pcis_bus.araddr),
    .s_axi_arlen   (sh_cl_dma_pcis_bus.arlen), 
    .s_axi_arvalid (sh_cl_dma_pcis_bus.arvalid),
    .s_axi_arsize  (sh_cl_dma_pcis_bus.arsize),
    .s_axi_arready (sh_cl_dma_pcis_bus.arready),
    .s_axi_rid     (sh_cl_dma_pcis_bus.rid),
    .s_axi_rdata   (sh_cl_dma_pcis_bus.rdata),
    .s_axi_rresp   (sh_cl_dma_pcis_bus.rresp),
    .s_axi_rlast   (sh_cl_dma_pcis_bus.rlast),
    .s_axi_rvalid  (sh_cl_dma_pcis_bus.rvalid),
    .s_axi_rready  (sh_cl_dma_pcis_bus.rready),

    .m_axi_awid    (sh_cl_dma_pcis_q.awid),
    .m_axi_awaddr  (sh_cl_dma_pcis_q.awaddr), 
    .m_axi_awlen   (sh_cl_dma_pcis_q.awlen),
    .m_axi_awvalid (sh_cl_dma_pcis_q.awvalid),
    .m_axi_awsize  (sh_cl_dma_pcis_q.awsize),
    .m_axi_awready (sh_cl_dma_pcis_q.awready),
    .m_axi_wdata   (sh_cl_dma_pcis_q.wdata),  
    .m_axi_wstrb   (sh_cl_dma_pcis_q.wstrb),
    .m_axi_wvalid  (sh_cl_dma_pcis_q.wvalid), 
    .m_axi_wlast   (sh_cl_dma_pcis_q.wlast),
    .m_axi_wready  (sh_cl_dma_pcis_q.wready), 
    .m_axi_bresp   (sh_cl_dma_pcis_q.bresp),  
    .m_axi_bvalid  (sh_cl_dma_pcis_q.bvalid), 
    .m_axi_bid     (sh_cl_dma_pcis_q.bid),
    .m_axi_bready  (sh_cl_dma_pcis_q.bready), 
    .m_axi_arid    (sh_cl_dma_pcis_q.arid), 
    .m_axi_araddr  (sh_cl_dma_pcis_q.araddr), 
    .m_axi_arlen   (sh_cl_dma_pcis_q.arlen), 
    .m_axi_arsize  (sh_cl_dma_pcis_q.arsize), 
    .m_axi_arvalid (sh_cl_dma_pcis_q.arvalid),
    .m_axi_arready (sh_cl_dma_pcis_q.arready),
    .m_axi_rid     (sh_cl_dma_pcis_q.rid),  
    .m_axi_rdata   (sh_cl_dma_pcis_q.rdata),  
    .m_axi_rresp   (sh_cl_dma_pcis_q.rresp),  
    .m_axi_rlast   (sh_cl_dma_pcis_q.rlast),  
    .m_axi_rvalid  (sh_cl_dma_pcis_q.rvalid), 
    .m_axi_rready  (sh_cl_dma_pcis_q.rready)
);

logic network_valid;
logic network_ready;
logic ar_sent = 0;
logic aw_sent = 0;
// fpga_pci_poke64
// fpga_pci_write_burst
sorter sort(
  .clock(clk_main_a0),
  .reset(!rst_main_n_sync),
  .io_blockValid(sh_cl_dma_pcis_wvalid && aw_sent),
  .io_block(sh_cl_dma_pcis_wdata),
  .io_downstreamReady(sh_cl_dma_pcis_rready && ar_sent),
  .io_thisReady(network_ready),
  .io_outValid(network_valid),
  .io_out(cl_sh_dma_pcis_rdata)
);

/*
always_ff @(posedge clk_main_a0) begin
  if (cl_sh_dma_pcis_wready && sh_cl_dma_pcis_wvalid) begin
    $display ("InData 0x%x...", sh_cl_dma_pcis_wdata);
  end
  if (sh_cl_dma_pcis_arvalid && cl_sh_dma_pcis_arready) begin
    $display ("Read address size/len 0x%x/0x%x...", sh_cl_dma_pcis_arsize, sh_cl_dma_pcis_arlen);
    $display ("Read address request 0x%x...", sh_cl_dma_pcis_araddr);
  end
  if (sh_cl_dma_pcis_awvalid && cl_sh_dma_pcis_awready) begin
    $display ("Write address 0x%x...", sh_cl_dma_pcis_awaddr);
  end
  if (sh_cl_dma_pcis_rready && cl_sh_dma_pcis_rvalid) begin
    $display ("OutData 0x%x...", cl_sh_dma_pcis_rdata);
    $display ("rlast 0x%x...", cl_sh_dma_pcis_rlast);
  end
  if (cl_sh_dma_pcis_bvalid && sh_cl_dma_pcis_bready) begin
    $display ("bvalid...");
  end
  if (sh_cl_dma_pcis_awvalid && cl_sh_dma_pcis_awready) begin
    $display ("aw_sent...");
  end
end
*/

// assign sh_cl_dma_pcis_bus.awvalid = sh_cl_dma_pcis_awvalid;
// assign sh_cl_dma_pcis_bus.awaddr = sh_cl_dma_pcis_awaddr;
// assign sh_cl_dma_pcis_bus.awid[5:0] = sh_cl_dma_pcis_awid;
// assign sh_cl_dma_pcis_bus.awlen = sh_cl_dma_pcis_awlen;
// assign sh_cl_dma_pcis_bus.awsize = sh_cl_dma_pcis_awsize;
// assign sh_cl_dma_pcis_bus.wvalid = sh_cl_dma_pcis_wvalid;
// assign sh_cl_dma_pcis_bus.wdata = sh_cl_dma_pcis_wdata;
// assign sh_cl_dma_pcis_bus.wstrb = sh_cl_dma_pcis_wstrb;
// assign sh_cl_dma_pcis_bus.wlast = sh_cl_dma_pcis_wlast;
// assign cl_sh_dma_pcis_wready = sh_cl_dma_pcis_bus.wready;
assign cl_sh_dma_pcis_bresp = 0;
// assign sh_cl_dma_pcis_bus.bready = sh_cl_dma_pcis_bready;
assign cl_sh_dma_pcis_bid = 0;
// assign sh_cl_dma_pcis_bus.arvalid = sh_cl_dma_pcis_arvalid;
// assign sh_cl_dma_pcis_bus.araddr = sh_cl_dma_pcis_araddr;
// assign sh_cl_dma_pcis_bus.arid[5:0] = sh_cl_dma_pcis_arid;
// assign sh_cl_dma_pcis_bus.arlen = sh_cl_dma_pcis_arlen;
// assign sh_cl_dma_pcis_bus.arsize = sh_cl_dma_pcis_arsize;
// assign cl_sh_dma_pcis_rvalid = sh_cl_dma_pcis_bus.rvalid;
assign cl_sh_dma_pcis_rid = 0;
assign cl_sh_dma_pcis_rresp = 0;
// assign cl_sh_dma_pcis_rdata = sh_cl_dma_pcis_bus.rdata;
// assign sh_cl_dma_pcis_bus.rready = sh_cl_dma_pcis_rready;

assign cl_sh_flr_done = 1;

logic [7:0] beat_count;
logic [7:0] arlen;
assign cl_sh_dma_pcis_arready = ar_sent == 0;
assign cl_sh_dma_pcis_rlast = beat_count == arlen;
assign cl_sh_dma_pcis_rvalid = ar_sent && network_valid;
always_ff @(posedge clk_main_a0) begin
  if (!rst_main_n_sync) begin
    ar_sent <= 0; 
  end
  else if (sh_cl_dma_pcis_arvalid && cl_sh_dma_pcis_arready) begin
    beat_count <= 0;
    arlen <= sh_cl_dma_pcis_arlen;
    ar_sent <= 1;
  end
  else if (sh_cl_dma_pcis_rready && cl_sh_dma_pcis_rvalid) begin
    if (cl_sh_dma_pcis_rlast) begin    
      ar_sent <= 0; 
    end
    else begin
      beat_count <= beat_count + 1;
    end
  end
end

logic bvalid = 0;
assign cl_sh_dma_pcis_awready = aw_sent == 0;
assign cl_sh_dma_pcis_wready = aw_sent && network_ready;
assign cl_sh_dma_pcis_bvalid = bvalid;
always_ff @(posedge clk_main_a0) begin
  if (!rst_main_n_sync) begin
    aw_sent <= 0; 
  end
  else if (sh_cl_dma_pcis_awvalid && cl_sh_dma_pcis_awready) begin
    aw_sent <= 1;
  end
  else if (bvalid && sh_cl_dma_pcis_bready) begin
    aw_sent <= 0;
  end
  bvalid <= bvalid && sh_cl_dma_pcis_bready
            ? 1'b0  : 
            ~bvalid && cl_sh_dma_pcis_wready && sh_cl_dma_pcis_wvalid && sh_cl_dma_pcis_wlast
            ? 1'b1  :
            bvalid;
end

/*
//-------------------------------------------------
// Hello World Register
//-------------------------------------------------
// When read it, returns the byte-flipped value.

always_ff @(posedge clk_main_a0)
   if (!rst_main_n_sync) begin                    // Reset
      hello_world_q[31:0] <= 32'h0000_0000;
   end
   else if (wready & (wr_addr == `HELLO_WORLD_REG_ADDR)) begin  
      hello_world_q[31:0] <= wdata[31:0];
   end
   else begin                                // Hold Value
      hello_world_q[31:0] <= hello_world_q[31:0];
   end

assign hello_world_q_byte_swapped[31:0] = {hello_world_q[7:0],   hello_world_q[15:8],
                                           hello_world_q[23:16], hello_world_q[31:24]};
*/

//-------------------------------------------------
// Virtual LED Register
//-------------------------------------------------
// Flop/synchronize interface signals
always_ff @(posedge clk_main_a0)
   if (!rst_main_n_sync) begin                    // Reset
      sh_cl_status_vdip_q[15:0]  <= 16'h0000;
      sh_cl_status_vdip_q2[15:0] <= 16'h0000;
      cl_sh_status_vled[15:0]    <= 16'h0000;
   end
   else begin
      sh_cl_status_vdip_q[15:0]  <= sh_cl_status_vdip[15:0];
      sh_cl_status_vdip_q2[15:0] <= sh_cl_status_vdip_q[15:0];
      cl_sh_status_vled[15:0]    <= pre_cl_sh_status_vled[15:0];
   end

// The register contains 16 read-only bits corresponding to 16 LED's.
// For this example, the virtual LED register shadows the hello_world
// register.
// The same LED values can be read from the CL to Shell interface
// by using the linux FPGA tool: $ fpga-get-virtual-led -S 0

always_ff @(posedge clk_main_a0)
   if (!rst_main_n_sync) begin                    // Reset
      vled_q[15:0] <= 16'h0000;
   end
   else begin
      vled_q[15:0] <= hello_world_q[15:0];
   end

// The Virtual LED outputs will be masked with the Virtual DIP switches.
assign pre_cl_sh_status_vled[15:0] = vled_q[15:0] & sh_cl_status_vdip_q2[15:0];

//-------------------------------------------
// Tie-Off Global Signals
//-------------------------------------------
`ifndef CL_VERSION
   `define CL_VERSION 32'hee_ee_ee_00
`endif  


  assign cl_sh_status0[31:0] =  32'h0000_0FF0;
  assign cl_sh_status1[31:0] = `CL_VERSION;

//-----------------------------------------------
// Debug bridge, used if need chipscope
//-----------------------------------------------
`ifndef DISABLE_CHIPSCOPE_DEBUG

// Flop for timing global clock counter
logic[63:0] sh_cl_glcount0_q;

always_ff @(posedge clk_main_a0)
   if (!rst_main_n_sync)
      sh_cl_glcount0_q <= 0;
   else
      sh_cl_glcount0_q <= sh_cl_glcount0;


// Integrated Logic Analyzers (ILA)
   ila_0 CL_ILA_0 (
                   .clk    (clk_main_a0),
                   .probe0 (sh_ocl_awvalid_q),
                   .probe1 (sh_ocl_awaddr_q ),
                   .probe2 (ocl_sh_awready_q),
                   .probe3 (sh_ocl_arvalid_q),
                   .probe4 (sh_ocl_araddr_q ),
                   .probe5 (ocl_sh_arready_q)
                   );

   ila_0 CL_ILA_1 (
                   .clk    (clk_main_a0),
                   .probe0 (ocl_sh_bvalid_q),
                   .probe1 (sh_cl_glcount0_q),
                   .probe2 (sh_ocl_bready_q),
                   .probe3 (ocl_sh_rvalid_q),
                   .probe4 ({32'b0,ocl_sh_rdata_q[31:0]}),
                   .probe5 (sh_ocl_rready_q)
                   );

// Debug Bridge 
 cl_debug_bridge CL_DEBUG_BRIDGE (
      .clk(clk_main_a0),
      .S_BSCAN_VEC_drck(drck),
      .S_BSCAN_VEC_shift(shift),
      .S_BSCAN_VEC_tdi(tdi),
      .S_BSCAN_VEC_update(update),
      .S_BSCAN_VEC_sel(sel),
      .S_BSCAN_VEC_tdo(tdo),
      .S_BSCAN_VEC_tms(tms),
      .S_BSCAN_VEC_tck(tck),
      .S_BSCAN_VEC_runtest(runtest),
      .S_BSCAN_VEC_reset(reset),
      .S_BSCAN_VEC_capture(capture),
      .S_BSCAN_VEC_bscanid(bscanid)
   );

//-----------------------------------------------
// VIO Example - Needs Chipscope
//-----------------------------------------------
   // Counter running at 125MHz
   
   logic      vo_cnt_enable;
   logic      vo_cnt_load;
   logic      vo_cnt_clear;
   logic      vo_cnt_oneshot;
   logic [7:0]  vo_tick_value;
   logic [15:0] vo_cnt_load_value;
   logic [15:0] vo_cnt_watermark;

   logic      vo_cnt_enable_q = 0;
   logic      vo_cnt_load_q = 0;
   logic      vo_cnt_clear_q = 0;
   logic      vo_cnt_oneshot_q = 0;
   logic [7:0]  vo_tick_value_q = 0;
   logic [15:0] vo_cnt_load_value_q = 0;
   logic [15:0] vo_cnt_watermark_q = 0;

   logic        vi_tick;
   logic        vi_cnt_ge_watermark;
   logic [7:0]  vi_tick_cnt = 0;
   logic [15:0] vi_cnt = 0;
   
   // Tick counter and main counter
   always @(posedge clk_main_a0) begin

      vo_cnt_enable_q     <= vo_cnt_enable    ;
      vo_cnt_load_q       <= vo_cnt_load      ;
      vo_cnt_clear_q      <= vo_cnt_clear     ;
      vo_cnt_oneshot_q    <= vo_cnt_oneshot   ;
      vo_tick_value_q     <= vo_tick_value    ;
      vo_cnt_load_value_q <= vo_cnt_load_value;
      vo_cnt_watermark_q  <= vo_cnt_watermark ;

      vi_tick_cnt = vo_cnt_clear_q ? 0 :
                    ~vo_cnt_enable_q ? vi_tick_cnt :
                    (vi_tick_cnt >= vo_tick_value_q) ? 0 :
                    vi_tick_cnt + 1;

      vi_cnt = vo_cnt_clear_q ? 0 :
               vo_cnt_load_q ? vo_cnt_load_value_q :
               ~vo_cnt_enable_q ? vi_cnt :
               (vi_tick_cnt >= vo_tick_value_q) && (~vo_cnt_oneshot_q || (vi_cnt <= 16'hFFFF)) ? vi_cnt + 1 :
               vi_cnt;

      vi_tick = (vi_tick_cnt >= vo_tick_value_q);

      vi_cnt_ge_watermark = (vi_cnt >= vo_cnt_watermark_q);
      
   end // always @ (posedge clk_main_a0)
   

   vio_0 CL_VIO_0 (
                   .clk    (clk_main_a0),
                   .probe_in0  (vi_tick),
                   .probe_in1  (vi_cnt_ge_watermark),
                   .probe_in2  (vi_tick_cnt),
                   .probe_in3  (vi_cnt),
                   .probe_out0 (vo_cnt_enable),
                   .probe_out1 (vo_cnt_load),
                   .probe_out2 (vo_cnt_clear),
                   .probe_out3 (vo_cnt_oneshot),
                   .probe_out4 (vo_tick_value),
                   .probe_out5 (vo_cnt_load_value),
                   .probe_out6 (vo_cnt_watermark)
                   );
   
   ila_vio_counter CL_VIO_ILA (
                   .clk     (clk_main_a0),
                   .probe0  (vi_tick),
                   .probe1  (vi_cnt_ge_watermark),
                   .probe2  (vi_tick_cnt),
                   .probe3  (vi_cnt),
                   .probe4  (vo_cnt_enable_q),
                   .probe5  (vo_cnt_load_q),
                   .probe6  (vo_cnt_clear_q),
                   .probe7  (vo_cnt_oneshot_q),
                   .probe8  (vo_tick_value_q),
                   .probe9  (vo_cnt_load_value_q),
                   .probe10 (vo_cnt_watermark_q)
                   );
   
`endif //  `ifndef DISABLE_CHIPSCOPE_DEBUG

endmodule





