`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module PassThrough(
  input   clock,
  input   reset,
  input  [511:0] io_inputMemBlock,
  input   io_inputMemBlockValid,
  input  [9:0] io_inputBits,
  output  io_inputMemConsumed,
  input   io_inputFinished,
  output [511:0] io_outputMemBlock,
  output  io_outputMemBlockValid,
  output [9:0] io_outputBits,
  output  io_outputFinished,
  input   io_outputMemFlushed
);
  reg  inputMemBlock_0;
  reg [31:0] _GEN_1539;
  reg  inputMemBlock_1;
  reg [31:0] _GEN_1540;
  reg  inputMemBlock_2;
  reg [31:0] _GEN_1541;
  reg  inputMemBlock_3;
  reg [31:0] _GEN_1542;
  reg  inputMemBlock_4;
  reg [31:0] _GEN_1543;
  reg  inputMemBlock_5;
  reg [31:0] _GEN_1544;
  reg  inputMemBlock_6;
  reg [31:0] _GEN_1545;
  reg  inputMemBlock_7;
  reg [31:0] _GEN_1546;
  reg  inputMemBlock_8;
  reg [31:0] _GEN_1547;
  reg  inputMemBlock_9;
  reg [31:0] _GEN_1548;
  reg  inputMemBlock_10;
  reg [31:0] _GEN_1549;
  reg  inputMemBlock_11;
  reg [31:0] _GEN_1550;
  reg  inputMemBlock_12;
  reg [31:0] _GEN_1551;
  reg  inputMemBlock_13;
  reg [31:0] _GEN_1552;
  reg  inputMemBlock_14;
  reg [31:0] _GEN_1553;
  reg  inputMemBlock_15;
  reg [31:0] _GEN_1554;
  reg  inputMemBlock_16;
  reg [31:0] _GEN_1555;
  reg  inputMemBlock_17;
  reg [31:0] _GEN_1556;
  reg  inputMemBlock_18;
  reg [31:0] _GEN_1557;
  reg  inputMemBlock_19;
  reg [31:0] _GEN_1558;
  reg  inputMemBlock_20;
  reg [31:0] _GEN_1559;
  reg  inputMemBlock_21;
  reg [31:0] _GEN_1560;
  reg  inputMemBlock_22;
  reg [31:0] _GEN_1561;
  reg  inputMemBlock_23;
  reg [31:0] _GEN_1562;
  reg  inputMemBlock_24;
  reg [31:0] _GEN_1563;
  reg  inputMemBlock_25;
  reg [31:0] _GEN_1564;
  reg  inputMemBlock_26;
  reg [31:0] _GEN_1565;
  reg  inputMemBlock_27;
  reg [31:0] _GEN_1566;
  reg  inputMemBlock_28;
  reg [31:0] _GEN_1567;
  reg  inputMemBlock_29;
  reg [31:0] _GEN_1568;
  reg  inputMemBlock_30;
  reg [31:0] _GEN_1569;
  reg  inputMemBlock_31;
  reg [31:0] _GEN_1570;
  reg  inputMemBlock_32;
  reg [31:0] _GEN_1571;
  reg  inputMemBlock_33;
  reg [31:0] _GEN_1572;
  reg  inputMemBlock_34;
  reg [31:0] _GEN_1573;
  reg  inputMemBlock_35;
  reg [31:0] _GEN_1574;
  reg  inputMemBlock_36;
  reg [31:0] _GEN_1575;
  reg  inputMemBlock_37;
  reg [31:0] _GEN_1576;
  reg  inputMemBlock_38;
  reg [31:0] _GEN_1577;
  reg  inputMemBlock_39;
  reg [31:0] _GEN_1578;
  reg  inputMemBlock_40;
  reg [31:0] _GEN_1579;
  reg  inputMemBlock_41;
  reg [31:0] _GEN_1580;
  reg  inputMemBlock_42;
  reg [31:0] _GEN_1581;
  reg  inputMemBlock_43;
  reg [31:0] _GEN_1582;
  reg  inputMemBlock_44;
  reg [31:0] _GEN_1583;
  reg  inputMemBlock_45;
  reg [31:0] _GEN_1584;
  reg  inputMemBlock_46;
  reg [31:0] _GEN_1585;
  reg  inputMemBlock_47;
  reg [31:0] _GEN_1586;
  reg  inputMemBlock_48;
  reg [31:0] _GEN_1587;
  reg  inputMemBlock_49;
  reg [31:0] _GEN_1588;
  reg  inputMemBlock_50;
  reg [31:0] _GEN_1589;
  reg  inputMemBlock_51;
  reg [31:0] _GEN_1590;
  reg  inputMemBlock_52;
  reg [31:0] _GEN_1591;
  reg  inputMemBlock_53;
  reg [31:0] _GEN_1592;
  reg  inputMemBlock_54;
  reg [31:0] _GEN_1593;
  reg  inputMemBlock_55;
  reg [31:0] _GEN_1594;
  reg  inputMemBlock_56;
  reg [31:0] _GEN_1595;
  reg  inputMemBlock_57;
  reg [31:0] _GEN_1596;
  reg  inputMemBlock_58;
  reg [31:0] _GEN_1597;
  reg  inputMemBlock_59;
  reg [31:0] _GEN_1598;
  reg  inputMemBlock_60;
  reg [31:0] _GEN_1599;
  reg  inputMemBlock_61;
  reg [31:0] _GEN_1600;
  reg  inputMemBlock_62;
  reg [31:0] _GEN_1601;
  reg  inputMemBlock_63;
  reg [31:0] _GEN_1602;
  reg  inputMemBlock_64;
  reg [31:0] _GEN_1603;
  reg  inputMemBlock_65;
  reg [31:0] _GEN_1604;
  reg  inputMemBlock_66;
  reg [31:0] _GEN_1605;
  reg  inputMemBlock_67;
  reg [31:0] _GEN_1606;
  reg  inputMemBlock_68;
  reg [31:0] _GEN_1607;
  reg  inputMemBlock_69;
  reg [31:0] _GEN_1608;
  reg  inputMemBlock_70;
  reg [31:0] _GEN_1609;
  reg  inputMemBlock_71;
  reg [31:0] _GEN_1610;
  reg  inputMemBlock_72;
  reg [31:0] _GEN_1611;
  reg  inputMemBlock_73;
  reg [31:0] _GEN_1612;
  reg  inputMemBlock_74;
  reg [31:0] _GEN_1613;
  reg  inputMemBlock_75;
  reg [31:0] _GEN_1614;
  reg  inputMemBlock_76;
  reg [31:0] _GEN_1615;
  reg  inputMemBlock_77;
  reg [31:0] _GEN_1616;
  reg  inputMemBlock_78;
  reg [31:0] _GEN_1617;
  reg  inputMemBlock_79;
  reg [31:0] _GEN_1618;
  reg  inputMemBlock_80;
  reg [31:0] _GEN_1619;
  reg  inputMemBlock_81;
  reg [31:0] _GEN_1620;
  reg  inputMemBlock_82;
  reg [31:0] _GEN_1621;
  reg  inputMemBlock_83;
  reg [31:0] _GEN_1622;
  reg  inputMemBlock_84;
  reg [31:0] _GEN_1623;
  reg  inputMemBlock_85;
  reg [31:0] _GEN_1624;
  reg  inputMemBlock_86;
  reg [31:0] _GEN_1625;
  reg  inputMemBlock_87;
  reg [31:0] _GEN_1626;
  reg  inputMemBlock_88;
  reg [31:0] _GEN_1627;
  reg  inputMemBlock_89;
  reg [31:0] _GEN_1628;
  reg  inputMemBlock_90;
  reg [31:0] _GEN_1629;
  reg  inputMemBlock_91;
  reg [31:0] _GEN_1630;
  reg  inputMemBlock_92;
  reg [31:0] _GEN_1631;
  reg  inputMemBlock_93;
  reg [31:0] _GEN_1632;
  reg  inputMemBlock_94;
  reg [31:0] _GEN_1633;
  reg  inputMemBlock_95;
  reg [31:0] _GEN_1634;
  reg  inputMemBlock_96;
  reg [31:0] _GEN_1635;
  reg  inputMemBlock_97;
  reg [31:0] _GEN_1636;
  reg  inputMemBlock_98;
  reg [31:0] _GEN_1637;
  reg  inputMemBlock_99;
  reg [31:0] _GEN_1638;
  reg  inputMemBlock_100;
  reg [31:0] _GEN_1639;
  reg  inputMemBlock_101;
  reg [31:0] _GEN_1640;
  reg  inputMemBlock_102;
  reg [31:0] _GEN_1641;
  reg  inputMemBlock_103;
  reg [31:0] _GEN_1642;
  reg  inputMemBlock_104;
  reg [31:0] _GEN_1643;
  reg  inputMemBlock_105;
  reg [31:0] _GEN_1644;
  reg  inputMemBlock_106;
  reg [31:0] _GEN_1645;
  reg  inputMemBlock_107;
  reg [31:0] _GEN_1646;
  reg  inputMemBlock_108;
  reg [31:0] _GEN_1647;
  reg  inputMemBlock_109;
  reg [31:0] _GEN_1648;
  reg  inputMemBlock_110;
  reg [31:0] _GEN_1649;
  reg  inputMemBlock_111;
  reg [31:0] _GEN_1650;
  reg  inputMemBlock_112;
  reg [31:0] _GEN_1651;
  reg  inputMemBlock_113;
  reg [31:0] _GEN_1652;
  reg  inputMemBlock_114;
  reg [31:0] _GEN_1653;
  reg  inputMemBlock_115;
  reg [31:0] _GEN_1654;
  reg  inputMemBlock_116;
  reg [31:0] _GEN_1655;
  reg  inputMemBlock_117;
  reg [31:0] _GEN_1656;
  reg  inputMemBlock_118;
  reg [31:0] _GEN_1657;
  reg  inputMemBlock_119;
  reg [31:0] _GEN_1658;
  reg  inputMemBlock_120;
  reg [31:0] _GEN_1659;
  reg  inputMemBlock_121;
  reg [31:0] _GEN_1660;
  reg  inputMemBlock_122;
  reg [31:0] _GEN_1661;
  reg  inputMemBlock_123;
  reg [31:0] _GEN_1662;
  reg  inputMemBlock_124;
  reg [31:0] _GEN_1663;
  reg  inputMemBlock_125;
  reg [31:0] _GEN_1664;
  reg  inputMemBlock_126;
  reg [31:0] _GEN_1665;
  reg  inputMemBlock_127;
  reg [31:0] _GEN_1666;
  reg  inputMemBlock_128;
  reg [31:0] _GEN_1667;
  reg  inputMemBlock_129;
  reg [31:0] _GEN_1668;
  reg  inputMemBlock_130;
  reg [31:0] _GEN_1669;
  reg  inputMemBlock_131;
  reg [31:0] _GEN_1670;
  reg  inputMemBlock_132;
  reg [31:0] _GEN_1671;
  reg  inputMemBlock_133;
  reg [31:0] _GEN_1672;
  reg  inputMemBlock_134;
  reg [31:0] _GEN_1673;
  reg  inputMemBlock_135;
  reg [31:0] _GEN_1674;
  reg  inputMemBlock_136;
  reg [31:0] _GEN_1675;
  reg  inputMemBlock_137;
  reg [31:0] _GEN_1676;
  reg  inputMemBlock_138;
  reg [31:0] _GEN_1677;
  reg  inputMemBlock_139;
  reg [31:0] _GEN_1678;
  reg  inputMemBlock_140;
  reg [31:0] _GEN_1679;
  reg  inputMemBlock_141;
  reg [31:0] _GEN_1680;
  reg  inputMemBlock_142;
  reg [31:0] _GEN_1681;
  reg  inputMemBlock_143;
  reg [31:0] _GEN_1682;
  reg  inputMemBlock_144;
  reg [31:0] _GEN_1683;
  reg  inputMemBlock_145;
  reg [31:0] _GEN_1684;
  reg  inputMemBlock_146;
  reg [31:0] _GEN_1685;
  reg  inputMemBlock_147;
  reg [31:0] _GEN_1686;
  reg  inputMemBlock_148;
  reg [31:0] _GEN_1687;
  reg  inputMemBlock_149;
  reg [31:0] _GEN_1688;
  reg  inputMemBlock_150;
  reg [31:0] _GEN_1689;
  reg  inputMemBlock_151;
  reg [31:0] _GEN_1690;
  reg  inputMemBlock_152;
  reg [31:0] _GEN_1691;
  reg  inputMemBlock_153;
  reg [31:0] _GEN_1692;
  reg  inputMemBlock_154;
  reg [31:0] _GEN_1693;
  reg  inputMemBlock_155;
  reg [31:0] _GEN_1694;
  reg  inputMemBlock_156;
  reg [31:0] _GEN_1695;
  reg  inputMemBlock_157;
  reg [31:0] _GEN_1696;
  reg  inputMemBlock_158;
  reg [31:0] _GEN_1697;
  reg  inputMemBlock_159;
  reg [31:0] _GEN_1698;
  reg  inputMemBlock_160;
  reg [31:0] _GEN_1699;
  reg  inputMemBlock_161;
  reg [31:0] _GEN_1700;
  reg  inputMemBlock_162;
  reg [31:0] _GEN_1701;
  reg  inputMemBlock_163;
  reg [31:0] _GEN_1702;
  reg  inputMemBlock_164;
  reg [31:0] _GEN_1703;
  reg  inputMemBlock_165;
  reg [31:0] _GEN_1704;
  reg  inputMemBlock_166;
  reg [31:0] _GEN_1705;
  reg  inputMemBlock_167;
  reg [31:0] _GEN_1706;
  reg  inputMemBlock_168;
  reg [31:0] _GEN_1707;
  reg  inputMemBlock_169;
  reg [31:0] _GEN_1708;
  reg  inputMemBlock_170;
  reg [31:0] _GEN_1709;
  reg  inputMemBlock_171;
  reg [31:0] _GEN_1710;
  reg  inputMemBlock_172;
  reg [31:0] _GEN_1711;
  reg  inputMemBlock_173;
  reg [31:0] _GEN_1712;
  reg  inputMemBlock_174;
  reg [31:0] _GEN_1713;
  reg  inputMemBlock_175;
  reg [31:0] _GEN_1714;
  reg  inputMemBlock_176;
  reg [31:0] _GEN_1715;
  reg  inputMemBlock_177;
  reg [31:0] _GEN_1716;
  reg  inputMemBlock_178;
  reg [31:0] _GEN_1717;
  reg  inputMemBlock_179;
  reg [31:0] _GEN_1718;
  reg  inputMemBlock_180;
  reg [31:0] _GEN_1719;
  reg  inputMemBlock_181;
  reg [31:0] _GEN_1720;
  reg  inputMemBlock_182;
  reg [31:0] _GEN_1721;
  reg  inputMemBlock_183;
  reg [31:0] _GEN_1722;
  reg  inputMemBlock_184;
  reg [31:0] _GEN_1723;
  reg  inputMemBlock_185;
  reg [31:0] _GEN_1724;
  reg  inputMemBlock_186;
  reg [31:0] _GEN_1725;
  reg  inputMemBlock_187;
  reg [31:0] _GEN_1726;
  reg  inputMemBlock_188;
  reg [31:0] _GEN_1727;
  reg  inputMemBlock_189;
  reg [31:0] _GEN_1728;
  reg  inputMemBlock_190;
  reg [31:0] _GEN_1729;
  reg  inputMemBlock_191;
  reg [31:0] _GEN_1730;
  reg  inputMemBlock_192;
  reg [31:0] _GEN_1731;
  reg  inputMemBlock_193;
  reg [31:0] _GEN_1732;
  reg  inputMemBlock_194;
  reg [31:0] _GEN_1733;
  reg  inputMemBlock_195;
  reg [31:0] _GEN_1734;
  reg  inputMemBlock_196;
  reg [31:0] _GEN_1735;
  reg  inputMemBlock_197;
  reg [31:0] _GEN_1736;
  reg  inputMemBlock_198;
  reg [31:0] _GEN_1737;
  reg  inputMemBlock_199;
  reg [31:0] _GEN_1738;
  reg  inputMemBlock_200;
  reg [31:0] _GEN_1739;
  reg  inputMemBlock_201;
  reg [31:0] _GEN_1740;
  reg  inputMemBlock_202;
  reg [31:0] _GEN_1741;
  reg  inputMemBlock_203;
  reg [31:0] _GEN_1742;
  reg  inputMemBlock_204;
  reg [31:0] _GEN_1743;
  reg  inputMemBlock_205;
  reg [31:0] _GEN_1744;
  reg  inputMemBlock_206;
  reg [31:0] _GEN_1745;
  reg  inputMemBlock_207;
  reg [31:0] _GEN_1746;
  reg  inputMemBlock_208;
  reg [31:0] _GEN_1747;
  reg  inputMemBlock_209;
  reg [31:0] _GEN_1748;
  reg  inputMemBlock_210;
  reg [31:0] _GEN_1749;
  reg  inputMemBlock_211;
  reg [31:0] _GEN_1750;
  reg  inputMemBlock_212;
  reg [31:0] _GEN_1751;
  reg  inputMemBlock_213;
  reg [31:0] _GEN_1752;
  reg  inputMemBlock_214;
  reg [31:0] _GEN_1753;
  reg  inputMemBlock_215;
  reg [31:0] _GEN_1754;
  reg  inputMemBlock_216;
  reg [31:0] _GEN_1755;
  reg  inputMemBlock_217;
  reg [31:0] _GEN_1756;
  reg  inputMemBlock_218;
  reg [31:0] _GEN_1757;
  reg  inputMemBlock_219;
  reg [31:0] _GEN_1758;
  reg  inputMemBlock_220;
  reg [31:0] _GEN_1759;
  reg  inputMemBlock_221;
  reg [31:0] _GEN_1760;
  reg  inputMemBlock_222;
  reg [31:0] _GEN_1761;
  reg  inputMemBlock_223;
  reg [31:0] _GEN_1762;
  reg  inputMemBlock_224;
  reg [31:0] _GEN_1763;
  reg  inputMemBlock_225;
  reg [31:0] _GEN_1764;
  reg  inputMemBlock_226;
  reg [31:0] _GEN_1765;
  reg  inputMemBlock_227;
  reg [31:0] _GEN_1766;
  reg  inputMemBlock_228;
  reg [31:0] _GEN_1767;
  reg  inputMemBlock_229;
  reg [31:0] _GEN_1768;
  reg  inputMemBlock_230;
  reg [31:0] _GEN_1769;
  reg  inputMemBlock_231;
  reg [31:0] _GEN_1770;
  reg  inputMemBlock_232;
  reg [31:0] _GEN_1771;
  reg  inputMemBlock_233;
  reg [31:0] _GEN_1772;
  reg  inputMemBlock_234;
  reg [31:0] _GEN_1773;
  reg  inputMemBlock_235;
  reg [31:0] _GEN_1774;
  reg  inputMemBlock_236;
  reg [31:0] _GEN_1775;
  reg  inputMemBlock_237;
  reg [31:0] _GEN_1776;
  reg  inputMemBlock_238;
  reg [31:0] _GEN_1777;
  reg  inputMemBlock_239;
  reg [31:0] _GEN_1778;
  reg  inputMemBlock_240;
  reg [31:0] _GEN_1779;
  reg  inputMemBlock_241;
  reg [31:0] _GEN_1780;
  reg  inputMemBlock_242;
  reg [31:0] _GEN_1781;
  reg  inputMemBlock_243;
  reg [31:0] _GEN_1782;
  reg  inputMemBlock_244;
  reg [31:0] _GEN_1783;
  reg  inputMemBlock_245;
  reg [31:0] _GEN_1784;
  reg  inputMemBlock_246;
  reg [31:0] _GEN_1785;
  reg  inputMemBlock_247;
  reg [31:0] _GEN_1786;
  reg  inputMemBlock_248;
  reg [31:0] _GEN_1787;
  reg  inputMemBlock_249;
  reg [31:0] _GEN_1788;
  reg  inputMemBlock_250;
  reg [31:0] _GEN_1789;
  reg  inputMemBlock_251;
  reg [31:0] _GEN_1790;
  reg  inputMemBlock_252;
  reg [31:0] _GEN_1791;
  reg  inputMemBlock_253;
  reg [31:0] _GEN_1792;
  reg  inputMemBlock_254;
  reg [31:0] _GEN_1793;
  reg  inputMemBlock_255;
  reg [31:0] _GEN_1794;
  reg  inputMemBlock_256;
  reg [31:0] _GEN_1795;
  reg  inputMemBlock_257;
  reg [31:0] _GEN_1796;
  reg  inputMemBlock_258;
  reg [31:0] _GEN_1797;
  reg  inputMemBlock_259;
  reg [31:0] _GEN_1798;
  reg  inputMemBlock_260;
  reg [31:0] _GEN_1799;
  reg  inputMemBlock_261;
  reg [31:0] _GEN_1800;
  reg  inputMemBlock_262;
  reg [31:0] _GEN_1801;
  reg  inputMemBlock_263;
  reg [31:0] _GEN_1802;
  reg  inputMemBlock_264;
  reg [31:0] _GEN_1803;
  reg  inputMemBlock_265;
  reg [31:0] _GEN_1804;
  reg  inputMemBlock_266;
  reg [31:0] _GEN_1805;
  reg  inputMemBlock_267;
  reg [31:0] _GEN_1806;
  reg  inputMemBlock_268;
  reg [31:0] _GEN_1807;
  reg  inputMemBlock_269;
  reg [31:0] _GEN_1808;
  reg  inputMemBlock_270;
  reg [31:0] _GEN_1809;
  reg  inputMemBlock_271;
  reg [31:0] _GEN_1810;
  reg  inputMemBlock_272;
  reg [31:0] _GEN_1811;
  reg  inputMemBlock_273;
  reg [31:0] _GEN_1812;
  reg  inputMemBlock_274;
  reg [31:0] _GEN_1813;
  reg  inputMemBlock_275;
  reg [31:0] _GEN_1814;
  reg  inputMemBlock_276;
  reg [31:0] _GEN_1815;
  reg  inputMemBlock_277;
  reg [31:0] _GEN_1816;
  reg  inputMemBlock_278;
  reg [31:0] _GEN_1817;
  reg  inputMemBlock_279;
  reg [31:0] _GEN_1818;
  reg  inputMemBlock_280;
  reg [31:0] _GEN_1819;
  reg  inputMemBlock_281;
  reg [31:0] _GEN_1820;
  reg  inputMemBlock_282;
  reg [31:0] _GEN_1821;
  reg  inputMemBlock_283;
  reg [31:0] _GEN_1822;
  reg  inputMemBlock_284;
  reg [31:0] _GEN_1823;
  reg  inputMemBlock_285;
  reg [31:0] _GEN_1824;
  reg  inputMemBlock_286;
  reg [31:0] _GEN_1825;
  reg  inputMemBlock_287;
  reg [31:0] _GEN_1826;
  reg  inputMemBlock_288;
  reg [31:0] _GEN_1827;
  reg  inputMemBlock_289;
  reg [31:0] _GEN_1828;
  reg  inputMemBlock_290;
  reg [31:0] _GEN_1829;
  reg  inputMemBlock_291;
  reg [31:0] _GEN_1830;
  reg  inputMemBlock_292;
  reg [31:0] _GEN_1831;
  reg  inputMemBlock_293;
  reg [31:0] _GEN_1832;
  reg  inputMemBlock_294;
  reg [31:0] _GEN_1833;
  reg  inputMemBlock_295;
  reg [31:0] _GEN_1834;
  reg  inputMemBlock_296;
  reg [31:0] _GEN_1835;
  reg  inputMemBlock_297;
  reg [31:0] _GEN_1836;
  reg  inputMemBlock_298;
  reg [31:0] _GEN_1837;
  reg  inputMemBlock_299;
  reg [31:0] _GEN_1838;
  reg  inputMemBlock_300;
  reg [31:0] _GEN_1839;
  reg  inputMemBlock_301;
  reg [31:0] _GEN_1840;
  reg  inputMemBlock_302;
  reg [31:0] _GEN_1841;
  reg  inputMemBlock_303;
  reg [31:0] _GEN_1842;
  reg  inputMemBlock_304;
  reg [31:0] _GEN_1843;
  reg  inputMemBlock_305;
  reg [31:0] _GEN_1844;
  reg  inputMemBlock_306;
  reg [31:0] _GEN_1845;
  reg  inputMemBlock_307;
  reg [31:0] _GEN_1846;
  reg  inputMemBlock_308;
  reg [31:0] _GEN_1847;
  reg  inputMemBlock_309;
  reg [31:0] _GEN_1848;
  reg  inputMemBlock_310;
  reg [31:0] _GEN_1849;
  reg  inputMemBlock_311;
  reg [31:0] _GEN_1850;
  reg  inputMemBlock_312;
  reg [31:0] _GEN_1851;
  reg  inputMemBlock_313;
  reg [31:0] _GEN_1852;
  reg  inputMemBlock_314;
  reg [31:0] _GEN_1853;
  reg  inputMemBlock_315;
  reg [31:0] _GEN_1854;
  reg  inputMemBlock_316;
  reg [31:0] _GEN_1855;
  reg  inputMemBlock_317;
  reg [31:0] _GEN_1856;
  reg  inputMemBlock_318;
  reg [31:0] _GEN_1857;
  reg  inputMemBlock_319;
  reg [31:0] _GEN_1858;
  reg  inputMemBlock_320;
  reg [31:0] _GEN_1859;
  reg  inputMemBlock_321;
  reg [31:0] _GEN_1860;
  reg  inputMemBlock_322;
  reg [31:0] _GEN_1861;
  reg  inputMemBlock_323;
  reg [31:0] _GEN_1862;
  reg  inputMemBlock_324;
  reg [31:0] _GEN_1863;
  reg  inputMemBlock_325;
  reg [31:0] _GEN_1864;
  reg  inputMemBlock_326;
  reg [31:0] _GEN_1865;
  reg  inputMemBlock_327;
  reg [31:0] _GEN_1866;
  reg  inputMemBlock_328;
  reg [31:0] _GEN_1867;
  reg  inputMemBlock_329;
  reg [31:0] _GEN_1868;
  reg  inputMemBlock_330;
  reg [31:0] _GEN_1869;
  reg  inputMemBlock_331;
  reg [31:0] _GEN_1870;
  reg  inputMemBlock_332;
  reg [31:0] _GEN_1871;
  reg  inputMemBlock_333;
  reg [31:0] _GEN_1872;
  reg  inputMemBlock_334;
  reg [31:0] _GEN_1873;
  reg  inputMemBlock_335;
  reg [31:0] _GEN_1874;
  reg  inputMemBlock_336;
  reg [31:0] _GEN_1875;
  reg  inputMemBlock_337;
  reg [31:0] _GEN_1876;
  reg  inputMemBlock_338;
  reg [31:0] _GEN_1877;
  reg  inputMemBlock_339;
  reg [31:0] _GEN_1878;
  reg  inputMemBlock_340;
  reg [31:0] _GEN_1879;
  reg  inputMemBlock_341;
  reg [31:0] _GEN_1880;
  reg  inputMemBlock_342;
  reg [31:0] _GEN_1881;
  reg  inputMemBlock_343;
  reg [31:0] _GEN_1882;
  reg  inputMemBlock_344;
  reg [31:0] _GEN_1883;
  reg  inputMemBlock_345;
  reg [31:0] _GEN_1884;
  reg  inputMemBlock_346;
  reg [31:0] _GEN_1885;
  reg  inputMemBlock_347;
  reg [31:0] _GEN_1886;
  reg  inputMemBlock_348;
  reg [31:0] _GEN_1887;
  reg  inputMemBlock_349;
  reg [31:0] _GEN_1888;
  reg  inputMemBlock_350;
  reg [31:0] _GEN_1889;
  reg  inputMemBlock_351;
  reg [31:0] _GEN_1890;
  reg  inputMemBlock_352;
  reg [31:0] _GEN_1891;
  reg  inputMemBlock_353;
  reg [31:0] _GEN_1892;
  reg  inputMemBlock_354;
  reg [31:0] _GEN_1893;
  reg  inputMemBlock_355;
  reg [31:0] _GEN_1894;
  reg  inputMemBlock_356;
  reg [31:0] _GEN_1895;
  reg  inputMemBlock_357;
  reg [31:0] _GEN_1896;
  reg  inputMemBlock_358;
  reg [31:0] _GEN_1897;
  reg  inputMemBlock_359;
  reg [31:0] _GEN_1898;
  reg  inputMemBlock_360;
  reg [31:0] _GEN_1899;
  reg  inputMemBlock_361;
  reg [31:0] _GEN_1900;
  reg  inputMemBlock_362;
  reg [31:0] _GEN_1901;
  reg  inputMemBlock_363;
  reg [31:0] _GEN_1902;
  reg  inputMemBlock_364;
  reg [31:0] _GEN_1903;
  reg  inputMemBlock_365;
  reg [31:0] _GEN_1904;
  reg  inputMemBlock_366;
  reg [31:0] _GEN_1905;
  reg  inputMemBlock_367;
  reg [31:0] _GEN_1906;
  reg  inputMemBlock_368;
  reg [31:0] _GEN_1907;
  reg  inputMemBlock_369;
  reg [31:0] _GEN_1908;
  reg  inputMemBlock_370;
  reg [31:0] _GEN_1909;
  reg  inputMemBlock_371;
  reg [31:0] _GEN_1910;
  reg  inputMemBlock_372;
  reg [31:0] _GEN_1911;
  reg  inputMemBlock_373;
  reg [31:0] _GEN_1912;
  reg  inputMemBlock_374;
  reg [31:0] _GEN_1913;
  reg  inputMemBlock_375;
  reg [31:0] _GEN_1914;
  reg  inputMemBlock_376;
  reg [31:0] _GEN_1915;
  reg  inputMemBlock_377;
  reg [31:0] _GEN_1916;
  reg  inputMemBlock_378;
  reg [31:0] _GEN_1917;
  reg  inputMemBlock_379;
  reg [31:0] _GEN_1918;
  reg  inputMemBlock_380;
  reg [31:0] _GEN_1919;
  reg  inputMemBlock_381;
  reg [31:0] _GEN_1920;
  reg  inputMemBlock_382;
  reg [31:0] _GEN_1921;
  reg  inputMemBlock_383;
  reg [31:0] _GEN_1922;
  reg  inputMemBlock_384;
  reg [31:0] _GEN_1923;
  reg  inputMemBlock_385;
  reg [31:0] _GEN_1924;
  reg  inputMemBlock_386;
  reg [31:0] _GEN_1925;
  reg  inputMemBlock_387;
  reg [31:0] _GEN_1926;
  reg  inputMemBlock_388;
  reg [31:0] _GEN_1927;
  reg  inputMemBlock_389;
  reg [31:0] _GEN_1928;
  reg  inputMemBlock_390;
  reg [31:0] _GEN_1929;
  reg  inputMemBlock_391;
  reg [31:0] _GEN_1930;
  reg  inputMemBlock_392;
  reg [31:0] _GEN_1931;
  reg  inputMemBlock_393;
  reg [31:0] _GEN_1932;
  reg  inputMemBlock_394;
  reg [31:0] _GEN_1933;
  reg  inputMemBlock_395;
  reg [31:0] _GEN_1934;
  reg  inputMemBlock_396;
  reg [31:0] _GEN_1935;
  reg  inputMemBlock_397;
  reg [31:0] _GEN_1936;
  reg  inputMemBlock_398;
  reg [31:0] _GEN_1937;
  reg  inputMemBlock_399;
  reg [31:0] _GEN_1938;
  reg  inputMemBlock_400;
  reg [31:0] _GEN_1939;
  reg  inputMemBlock_401;
  reg [31:0] _GEN_1940;
  reg  inputMemBlock_402;
  reg [31:0] _GEN_1941;
  reg  inputMemBlock_403;
  reg [31:0] _GEN_1942;
  reg  inputMemBlock_404;
  reg [31:0] _GEN_1943;
  reg  inputMemBlock_405;
  reg [31:0] _GEN_1944;
  reg  inputMemBlock_406;
  reg [31:0] _GEN_1945;
  reg  inputMemBlock_407;
  reg [31:0] _GEN_1946;
  reg  inputMemBlock_408;
  reg [31:0] _GEN_1947;
  reg  inputMemBlock_409;
  reg [31:0] _GEN_1948;
  reg  inputMemBlock_410;
  reg [31:0] _GEN_1949;
  reg  inputMemBlock_411;
  reg [31:0] _GEN_1950;
  reg  inputMemBlock_412;
  reg [31:0] _GEN_1951;
  reg  inputMemBlock_413;
  reg [31:0] _GEN_1952;
  reg  inputMemBlock_414;
  reg [31:0] _GEN_1953;
  reg  inputMemBlock_415;
  reg [31:0] _GEN_1954;
  reg  inputMemBlock_416;
  reg [31:0] _GEN_1955;
  reg  inputMemBlock_417;
  reg [31:0] _GEN_1956;
  reg  inputMemBlock_418;
  reg [31:0] _GEN_1957;
  reg  inputMemBlock_419;
  reg [31:0] _GEN_1958;
  reg  inputMemBlock_420;
  reg [31:0] _GEN_1959;
  reg  inputMemBlock_421;
  reg [31:0] _GEN_1960;
  reg  inputMemBlock_422;
  reg [31:0] _GEN_1961;
  reg  inputMemBlock_423;
  reg [31:0] _GEN_1962;
  reg  inputMemBlock_424;
  reg [31:0] _GEN_1963;
  reg  inputMemBlock_425;
  reg [31:0] _GEN_1964;
  reg  inputMemBlock_426;
  reg [31:0] _GEN_1965;
  reg  inputMemBlock_427;
  reg [31:0] _GEN_1966;
  reg  inputMemBlock_428;
  reg [31:0] _GEN_1967;
  reg  inputMemBlock_429;
  reg [31:0] _GEN_1968;
  reg  inputMemBlock_430;
  reg [31:0] _GEN_1969;
  reg  inputMemBlock_431;
  reg [31:0] _GEN_1970;
  reg  inputMemBlock_432;
  reg [31:0] _GEN_1971;
  reg  inputMemBlock_433;
  reg [31:0] _GEN_1972;
  reg  inputMemBlock_434;
  reg [31:0] _GEN_1973;
  reg  inputMemBlock_435;
  reg [31:0] _GEN_1974;
  reg  inputMemBlock_436;
  reg [31:0] _GEN_1975;
  reg  inputMemBlock_437;
  reg [31:0] _GEN_1976;
  reg  inputMemBlock_438;
  reg [31:0] _GEN_1977;
  reg  inputMemBlock_439;
  reg [31:0] _GEN_1978;
  reg  inputMemBlock_440;
  reg [31:0] _GEN_1979;
  reg  inputMemBlock_441;
  reg [31:0] _GEN_1980;
  reg  inputMemBlock_442;
  reg [31:0] _GEN_1981;
  reg  inputMemBlock_443;
  reg [31:0] _GEN_1982;
  reg  inputMemBlock_444;
  reg [31:0] _GEN_1983;
  reg  inputMemBlock_445;
  reg [31:0] _GEN_1984;
  reg  inputMemBlock_446;
  reg [31:0] _GEN_1985;
  reg  inputMemBlock_447;
  reg [31:0] _GEN_1986;
  reg  inputMemBlock_448;
  reg [31:0] _GEN_1987;
  reg  inputMemBlock_449;
  reg [31:0] _GEN_1988;
  reg  inputMemBlock_450;
  reg [31:0] _GEN_1989;
  reg  inputMemBlock_451;
  reg [31:0] _GEN_1990;
  reg  inputMemBlock_452;
  reg [31:0] _GEN_1991;
  reg  inputMemBlock_453;
  reg [31:0] _GEN_1992;
  reg  inputMemBlock_454;
  reg [31:0] _GEN_1993;
  reg  inputMemBlock_455;
  reg [31:0] _GEN_1994;
  reg  inputMemBlock_456;
  reg [31:0] _GEN_1995;
  reg  inputMemBlock_457;
  reg [31:0] _GEN_1996;
  reg  inputMemBlock_458;
  reg [31:0] _GEN_1997;
  reg  inputMemBlock_459;
  reg [31:0] _GEN_1998;
  reg  inputMemBlock_460;
  reg [31:0] _GEN_1999;
  reg  inputMemBlock_461;
  reg [31:0] _GEN_2000;
  reg  inputMemBlock_462;
  reg [31:0] _GEN_2001;
  reg  inputMemBlock_463;
  reg [31:0] _GEN_2002;
  reg  inputMemBlock_464;
  reg [31:0] _GEN_2003;
  reg  inputMemBlock_465;
  reg [31:0] _GEN_2004;
  reg  inputMemBlock_466;
  reg [31:0] _GEN_2005;
  reg  inputMemBlock_467;
  reg [31:0] _GEN_2006;
  reg  inputMemBlock_468;
  reg [31:0] _GEN_2007;
  reg  inputMemBlock_469;
  reg [31:0] _GEN_2008;
  reg  inputMemBlock_470;
  reg [31:0] _GEN_2009;
  reg  inputMemBlock_471;
  reg [31:0] _GEN_2010;
  reg  inputMemBlock_472;
  reg [31:0] _GEN_2011;
  reg  inputMemBlock_473;
  reg [31:0] _GEN_2012;
  reg  inputMemBlock_474;
  reg [31:0] _GEN_2013;
  reg  inputMemBlock_475;
  reg [31:0] _GEN_2014;
  reg  inputMemBlock_476;
  reg [31:0] _GEN_2015;
  reg  inputMemBlock_477;
  reg [31:0] _GEN_2016;
  reg  inputMemBlock_478;
  reg [31:0] _GEN_2017;
  reg  inputMemBlock_479;
  reg [31:0] _GEN_2018;
  reg  inputMemBlock_480;
  reg [31:0] _GEN_2019;
  reg  inputMemBlock_481;
  reg [31:0] _GEN_2020;
  reg  inputMemBlock_482;
  reg [31:0] _GEN_2021;
  reg  inputMemBlock_483;
  reg [31:0] _GEN_2022;
  reg  inputMemBlock_484;
  reg [31:0] _GEN_2023;
  reg  inputMemBlock_485;
  reg [31:0] _GEN_2024;
  reg  inputMemBlock_486;
  reg [31:0] _GEN_2025;
  reg  inputMemBlock_487;
  reg [31:0] _GEN_2026;
  reg  inputMemBlock_488;
  reg [31:0] _GEN_2027;
  reg  inputMemBlock_489;
  reg [31:0] _GEN_2028;
  reg  inputMemBlock_490;
  reg [31:0] _GEN_2029;
  reg  inputMemBlock_491;
  reg [31:0] _GEN_2030;
  reg  inputMemBlock_492;
  reg [31:0] _GEN_2031;
  reg  inputMemBlock_493;
  reg [31:0] _GEN_2032;
  reg  inputMemBlock_494;
  reg [31:0] _GEN_2033;
  reg  inputMemBlock_495;
  reg [31:0] _GEN_2034;
  reg  inputMemBlock_496;
  reg [31:0] _GEN_2035;
  reg  inputMemBlock_497;
  reg [31:0] _GEN_2036;
  reg  inputMemBlock_498;
  reg [31:0] _GEN_2037;
  reg  inputMemBlock_499;
  reg [31:0] _GEN_2038;
  reg  inputMemBlock_500;
  reg [31:0] _GEN_2039;
  reg  inputMemBlock_501;
  reg [31:0] _GEN_2040;
  reg  inputMemBlock_502;
  reg [31:0] _GEN_2041;
  reg  inputMemBlock_503;
  reg [31:0] _GEN_2042;
  reg  inputMemBlock_504;
  reg [31:0] _GEN_2043;
  reg  inputMemBlock_505;
  reg [31:0] _GEN_2044;
  reg  inputMemBlock_506;
  reg [31:0] _GEN_2045;
  reg  inputMemBlock_507;
  reg [31:0] _GEN_2046;
  reg  inputMemBlock_508;
  reg [31:0] _GEN_2047;
  reg  inputMemBlock_509;
  reg [31:0] _GEN_2048;
  reg  inputMemBlock_510;
  reg [31:0] _GEN_2049;
  reg  inputMemBlock_511;
  reg [31:0] _GEN_2050;
  reg [9:0] inputBitsRemaining;
  reg [31:0] _GEN_2051;
  wire  _T_540;
  wire  _T_541;
  wire  _T_542;
  wire  _T_543;
  wire  _T_544;
  wire  _T_545;
  wire  _T_546;
  wire  _T_547;
  wire  _T_548;
  wire  _T_549;
  wire  _T_550;
  wire  _T_551;
  wire  _T_552;
  wire  _T_553;
  wire  _T_554;
  wire  _T_555;
  wire  _T_556;
  wire  _T_557;
  wire  _T_558;
  wire  _T_559;
  wire  _T_560;
  wire  _T_561;
  wire  _T_562;
  wire  _T_563;
  wire  _T_564;
  wire  _T_565;
  wire  _T_566;
  wire  _T_567;
  wire  _T_568;
  wire  _T_569;
  wire  _T_570;
  wire  _T_571;
  wire  _T_572;
  wire  _T_573;
  wire  _T_574;
  wire  _T_575;
  wire  _T_576;
  wire  _T_577;
  wire  _T_578;
  wire  _T_579;
  wire  _T_580;
  wire  _T_581;
  wire  _T_582;
  wire  _T_583;
  wire  _T_584;
  wire  _T_585;
  wire  _T_586;
  wire  _T_587;
  wire  _T_588;
  wire  _T_589;
  wire  _T_590;
  wire  _T_591;
  wire  _T_592;
  wire  _T_593;
  wire  _T_594;
  wire  _T_595;
  wire  _T_596;
  wire  _T_597;
  wire  _T_598;
  wire  _T_599;
  wire  _T_600;
  wire  _T_601;
  wire  _T_602;
  wire  _T_603;
  wire  _T_604;
  wire  _T_605;
  wire  _T_606;
  wire  _T_607;
  wire  _T_608;
  wire  _T_609;
  wire  _T_610;
  wire  _T_611;
  wire  _T_612;
  wire  _T_613;
  wire  _T_614;
  wire  _T_615;
  wire  _T_616;
  wire  _T_617;
  wire  _T_618;
  wire  _T_619;
  wire  _T_620;
  wire  _T_621;
  wire  _T_622;
  wire  _T_623;
  wire  _T_624;
  wire  _T_625;
  wire  _T_626;
  wire  _T_627;
  wire  _T_628;
  wire  _T_629;
  wire  _T_630;
  wire  _T_631;
  wire  _T_632;
  wire  _T_633;
  wire  _T_634;
  wire  _T_635;
  wire  _T_636;
  wire  _T_637;
  wire  _T_638;
  wire  _T_639;
  wire  _T_640;
  wire  _T_641;
  wire  _T_642;
  wire  _T_643;
  wire  _T_644;
  wire  _T_645;
  wire  _T_646;
  wire  _T_647;
  wire  _T_648;
  wire  _T_649;
  wire  _T_650;
  wire  _T_651;
  wire  _T_652;
  wire  _T_653;
  wire  _T_654;
  wire  _T_655;
  wire  _T_656;
  wire  _T_657;
  wire  _T_658;
  wire  _T_659;
  wire  _T_660;
  wire  _T_661;
  wire  _T_662;
  wire  _T_663;
  wire  _T_664;
  wire  _T_665;
  wire  _T_666;
  wire  _T_667;
  wire  _T_668;
  wire  _T_669;
  wire  _T_670;
  wire  _T_671;
  wire  _T_672;
  wire  _T_673;
  wire  _T_674;
  wire  _T_675;
  wire  _T_676;
  wire  _T_677;
  wire  _T_678;
  wire  _T_679;
  wire  _T_680;
  wire  _T_681;
  wire  _T_682;
  wire  _T_683;
  wire  _T_684;
  wire  _T_685;
  wire  _T_686;
  wire  _T_687;
  wire  _T_688;
  wire  _T_689;
  wire  _T_690;
  wire  _T_691;
  wire  _T_692;
  wire  _T_693;
  wire  _T_694;
  wire  _T_695;
  wire  _T_696;
  wire  _T_697;
  wire  _T_698;
  wire  _T_699;
  wire  _T_700;
  wire  _T_701;
  wire  _T_702;
  wire  _T_703;
  wire  _T_704;
  wire  _T_705;
  wire  _T_706;
  wire  _T_707;
  wire  _T_708;
  wire  _T_709;
  wire  _T_710;
  wire  _T_711;
  wire  _T_712;
  wire  _T_713;
  wire  _T_714;
  wire  _T_715;
  wire  _T_716;
  wire  _T_717;
  wire  _T_718;
  wire  _T_719;
  wire  _T_720;
  wire  _T_721;
  wire  _T_722;
  wire  _T_723;
  wire  _T_724;
  wire  _T_725;
  wire  _T_726;
  wire  _T_727;
  wire  _T_728;
  wire  _T_729;
  wire  _T_730;
  wire  _T_731;
  wire  _T_732;
  wire  _T_733;
  wire  _T_734;
  wire  _T_735;
  wire  _T_736;
  wire  _T_737;
  wire  _T_738;
  wire  _T_739;
  wire  _T_740;
  wire  _T_741;
  wire  _T_742;
  wire  _T_743;
  wire  _T_744;
  wire  _T_745;
  wire  _T_746;
  wire  _T_747;
  wire  _T_748;
  wire  _T_749;
  wire  _T_750;
  wire  _T_751;
  wire  _T_752;
  wire  _T_753;
  wire  _T_754;
  wire  _T_755;
  wire  _T_756;
  wire  _T_757;
  wire  _T_758;
  wire  _T_759;
  wire  _T_760;
  wire  _T_761;
  wire  _T_762;
  wire  _T_763;
  wire  _T_764;
  wire  _T_765;
  wire  _T_766;
  wire  _T_767;
  wire  _T_768;
  wire  _T_769;
  wire  _T_770;
  wire  _T_771;
  wire  _T_772;
  wire  _T_773;
  wire  _T_774;
  wire  _T_775;
  wire  _T_776;
  wire  _T_777;
  wire  _T_778;
  wire  _T_779;
  wire  _T_780;
  wire  _T_781;
  wire  _T_782;
  wire  _T_783;
  wire  _T_784;
  wire  _T_785;
  wire  _T_786;
  wire  _T_787;
  wire  _T_788;
  wire  _T_789;
  wire  _T_790;
  wire  _T_791;
  wire  _T_792;
  wire  _T_793;
  wire  _T_794;
  wire  _T_795;
  wire  _T_796;
  wire  _T_797;
  wire  _T_798;
  wire  _T_799;
  wire  _T_800;
  wire  _T_801;
  wire  _T_802;
  wire  _T_803;
  wire  _T_804;
  wire  _T_805;
  wire  _T_806;
  wire  _T_807;
  wire  _T_808;
  wire  _T_809;
  wire  _T_810;
  wire  _T_811;
  wire  _T_812;
  wire  _T_813;
  wire  _T_814;
  wire  _T_815;
  wire  _T_816;
  wire  _T_817;
  wire  _T_818;
  wire  _T_819;
  wire  _T_820;
  wire  _T_821;
  wire  _T_822;
  wire  _T_823;
  wire  _T_824;
  wire  _T_825;
  wire  _T_826;
  wire  _T_827;
  wire  _T_828;
  wire  _T_829;
  wire  _T_830;
  wire  _T_831;
  wire  _T_832;
  wire  _T_833;
  wire  _T_834;
  wire  _T_835;
  wire  _T_836;
  wire  _T_837;
  wire  _T_838;
  wire  _T_839;
  wire  _T_840;
  wire  _T_841;
  wire  _T_842;
  wire  _T_843;
  wire  _T_844;
  wire  _T_845;
  wire  _T_846;
  wire  _T_847;
  wire  _T_848;
  wire  _T_849;
  wire  _T_850;
  wire  _T_851;
  wire  _T_852;
  wire  _T_853;
  wire  _T_854;
  wire  _T_855;
  wire  _T_856;
  wire  _T_857;
  wire  _T_858;
  wire  _T_859;
  wire  _T_860;
  wire  _T_861;
  wire  _T_862;
  wire  _T_863;
  wire  _T_864;
  wire  _T_865;
  wire  _T_866;
  wire  _T_867;
  wire  _T_868;
  wire  _T_869;
  wire  _T_870;
  wire  _T_871;
  wire  _T_872;
  wire  _T_873;
  wire  _T_874;
  wire  _T_875;
  wire  _T_876;
  wire  _T_877;
  wire  _T_878;
  wire  _T_879;
  wire  _T_880;
  wire  _T_881;
  wire  _T_882;
  wire  _T_883;
  wire  _T_884;
  wire  _T_885;
  wire  _T_886;
  wire  _T_887;
  wire  _T_888;
  wire  _T_889;
  wire  _T_890;
  wire  _T_891;
  wire  _T_892;
  wire  _T_893;
  wire  _T_894;
  wire  _T_895;
  wire  _T_896;
  wire  _T_897;
  wire  _T_898;
  wire  _T_899;
  wire  _T_900;
  wire  _T_901;
  wire  _T_902;
  wire  _T_903;
  wire  _T_904;
  wire  _T_905;
  wire  _T_906;
  wire  _T_907;
  wire  _T_908;
  wire  _T_909;
  wire  _T_910;
  wire  _T_911;
  wire  _T_912;
  wire  _T_913;
  wire  _T_914;
  wire  _T_915;
  wire  _T_916;
  wire  _T_917;
  wire  _T_918;
  wire  _T_919;
  wire  _T_920;
  wire  _T_921;
  wire  _T_922;
  wire  _T_923;
  wire  _T_924;
  wire  _T_925;
  wire  _T_926;
  wire  _T_927;
  wire  _T_928;
  wire  _T_929;
  wire  _T_930;
  wire  _T_931;
  wire  _T_932;
  wire  _T_933;
  wire  _T_934;
  wire  _T_935;
  wire  _T_936;
  wire  _T_937;
  wire  _T_938;
  wire  _T_939;
  wire  _T_940;
  wire  _T_941;
  wire  _T_942;
  wire  _T_943;
  wire  _T_944;
  wire  _T_945;
  wire  _T_946;
  wire  _T_947;
  wire  _T_948;
  wire  _T_949;
  wire  _T_950;
  wire  _T_951;
  wire  _T_952;
  wire  _T_953;
  wire  _T_954;
  wire  _T_955;
  wire  _T_956;
  wire  _T_957;
  wire  _T_958;
  wire  _T_959;
  wire  _T_960;
  wire  _T_961;
  wire  _T_962;
  wire  _T_963;
  wire  _T_964;
  wire  _T_965;
  wire  _T_966;
  wire  _T_967;
  wire  _T_968;
  wire  _T_969;
  wire  _T_970;
  wire  _T_971;
  wire  _T_972;
  wire  _T_973;
  wire  _T_974;
  wire  _T_975;
  wire  _T_976;
  wire  _T_977;
  wire  _T_978;
  wire  _T_979;
  wire  _T_980;
  wire  _T_981;
  wire  _T_982;
  wire  _T_983;
  wire  _T_984;
  wire  _T_985;
  wire  _T_986;
  wire  _T_987;
  wire  _T_988;
  wire  _T_989;
  wire  _T_990;
  wire  _T_991;
  wire  _T_992;
  wire  _T_993;
  wire  _T_994;
  wire  _T_995;
  wire  _T_996;
  wire  _T_997;
  wire  _T_998;
  wire  _T_999;
  wire  _T_1000;
  wire  _T_1001;
  wire  _T_1002;
  wire  _T_1003;
  wire  _T_1004;
  wire  _T_1005;
  wire  _T_1006;
  wire  _T_1007;
  wire  _T_1008;
  wire  _T_1009;
  wire  _T_1010;
  wire  _T_1011;
  wire  _T_1012;
  wire  _T_1013;
  wire  _T_1014;
  wire  _T_1015;
  wire  _T_1016;
  wire  _T_1017;
  wire  _T_1018;
  wire  _T_1019;
  wire  _T_1020;
  wire  _T_1021;
  wire  _T_1022;
  wire  _T_1023;
  wire  _T_1024;
  wire  _T_1025;
  wire  _T_1026;
  wire  _T_1027;
  wire  _T_1028;
  wire  _T_1029;
  wire  _T_1030;
  wire  _T_1031;
  wire  _T_1032;
  wire  _T_1033;
  wire  _T_1034;
  wire  _T_1035;
  wire  _T_1036;
  wire  _T_1037;
  wire  _T_1038;
  wire  _T_1039;
  wire  _T_1040;
  wire  _T_1041;
  wire  _T_1042;
  wire  _T_1043;
  wire  _T_1044;
  wire  _T_1045;
  wire  _T_1046;
  wire  _T_1047;
  wire  _T_1048;
  wire  _T_1049;
  wire  _T_1050;
  wire  _T_1051;
  wire [9:0] _GEN_0;
  wire  _GEN_1;
  wire  _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire  _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire  _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_76;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire  _GEN_83;
  wire  _GEN_84;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire  _GEN_90;
  wire  _GEN_91;
  wire  _GEN_92;
  wire  _GEN_93;
  wire  _GEN_94;
  wire  _GEN_95;
  wire  _GEN_96;
  wire  _GEN_97;
  wire  _GEN_98;
  wire  _GEN_99;
  wire  _GEN_100;
  wire  _GEN_101;
  wire  _GEN_102;
  wire  _GEN_103;
  wire  _GEN_104;
  wire  _GEN_105;
  wire  _GEN_106;
  wire  _GEN_107;
  wire  _GEN_108;
  wire  _GEN_109;
  wire  _GEN_110;
  wire  _GEN_111;
  wire  _GEN_112;
  wire  _GEN_113;
  wire  _GEN_114;
  wire  _GEN_115;
  wire  _GEN_116;
  wire  _GEN_117;
  wire  _GEN_118;
  wire  _GEN_119;
  wire  _GEN_120;
  wire  _GEN_121;
  wire  _GEN_122;
  wire  _GEN_123;
  wire  _GEN_124;
  wire  _GEN_125;
  wire  _GEN_126;
  wire  _GEN_127;
  wire  _GEN_128;
  wire  _GEN_129;
  wire  _GEN_130;
  wire  _GEN_131;
  wire  _GEN_132;
  wire  _GEN_133;
  wire  _GEN_134;
  wire  _GEN_135;
  wire  _GEN_136;
  wire  _GEN_137;
  wire  _GEN_138;
  wire  _GEN_139;
  wire  _GEN_140;
  wire  _GEN_141;
  wire  _GEN_142;
  wire  _GEN_143;
  wire  _GEN_144;
  wire  _GEN_145;
  wire  _GEN_146;
  wire  _GEN_147;
  wire  _GEN_148;
  wire  _GEN_149;
  wire  _GEN_150;
  wire  _GEN_151;
  wire  _GEN_152;
  wire  _GEN_153;
  wire  _GEN_154;
  wire  _GEN_155;
  wire  _GEN_156;
  wire  _GEN_157;
  wire  _GEN_158;
  wire  _GEN_159;
  wire  _GEN_160;
  wire  _GEN_161;
  wire  _GEN_162;
  wire  _GEN_163;
  wire  _GEN_164;
  wire  _GEN_165;
  wire  _GEN_166;
  wire  _GEN_167;
  wire  _GEN_168;
  wire  _GEN_169;
  wire  _GEN_170;
  wire  _GEN_171;
  wire  _GEN_172;
  wire  _GEN_173;
  wire  _GEN_174;
  wire  _GEN_175;
  wire  _GEN_176;
  wire  _GEN_177;
  wire  _GEN_178;
  wire  _GEN_179;
  wire  _GEN_180;
  wire  _GEN_181;
  wire  _GEN_182;
  wire  _GEN_183;
  wire  _GEN_184;
  wire  _GEN_185;
  wire  _GEN_186;
  wire  _GEN_187;
  wire  _GEN_188;
  wire  _GEN_189;
  wire  _GEN_190;
  wire  _GEN_191;
  wire  _GEN_192;
  wire  _GEN_193;
  wire  _GEN_194;
  wire  _GEN_195;
  wire  _GEN_196;
  wire  _GEN_197;
  wire  _GEN_198;
  wire  _GEN_199;
  wire  _GEN_200;
  wire  _GEN_201;
  wire  _GEN_202;
  wire  _GEN_203;
  wire  _GEN_204;
  wire  _GEN_205;
  wire  _GEN_206;
  wire  _GEN_207;
  wire  _GEN_208;
  wire  _GEN_209;
  wire  _GEN_210;
  wire  _GEN_211;
  wire  _GEN_212;
  wire  _GEN_213;
  wire  _GEN_214;
  wire  _GEN_215;
  wire  _GEN_216;
  wire  _GEN_217;
  wire  _GEN_218;
  wire  _GEN_219;
  wire  _GEN_220;
  wire  _GEN_221;
  wire  _GEN_222;
  wire  _GEN_223;
  wire  _GEN_224;
  wire  _GEN_225;
  wire  _GEN_226;
  wire  _GEN_227;
  wire  _GEN_228;
  wire  _GEN_229;
  wire  _GEN_230;
  wire  _GEN_231;
  wire  _GEN_232;
  wire  _GEN_233;
  wire  _GEN_234;
  wire  _GEN_235;
  wire  _GEN_236;
  wire  _GEN_237;
  wire  _GEN_238;
  wire  _GEN_239;
  wire  _GEN_240;
  wire  _GEN_241;
  wire  _GEN_242;
  wire  _GEN_243;
  wire  _GEN_244;
  wire  _GEN_245;
  wire  _GEN_246;
  wire  _GEN_247;
  wire  _GEN_248;
  wire  _GEN_249;
  wire  _GEN_250;
  wire  _GEN_251;
  wire  _GEN_252;
  wire  _GEN_253;
  wire  _GEN_254;
  wire  _GEN_255;
  wire  _GEN_256;
  wire  _GEN_257;
  wire  _GEN_258;
  wire  _GEN_259;
  wire  _GEN_260;
  wire  _GEN_261;
  wire  _GEN_262;
  wire  _GEN_263;
  wire  _GEN_264;
  wire  _GEN_265;
  wire  _GEN_266;
  wire  _GEN_267;
  wire  _GEN_268;
  wire  _GEN_269;
  wire  _GEN_270;
  wire  _GEN_271;
  wire  _GEN_272;
  wire  _GEN_273;
  wire  _GEN_274;
  wire  _GEN_275;
  wire  _GEN_276;
  wire  _GEN_277;
  wire  _GEN_278;
  wire  _GEN_279;
  wire  _GEN_280;
  wire  _GEN_281;
  wire  _GEN_282;
  wire  _GEN_283;
  wire  _GEN_284;
  wire  _GEN_285;
  wire  _GEN_286;
  wire  _GEN_287;
  wire  _GEN_288;
  wire  _GEN_289;
  wire  _GEN_290;
  wire  _GEN_291;
  wire  _GEN_292;
  wire  _GEN_293;
  wire  _GEN_294;
  wire  _GEN_295;
  wire  _GEN_296;
  wire  _GEN_297;
  wire  _GEN_298;
  wire  _GEN_299;
  wire  _GEN_300;
  wire  _GEN_301;
  wire  _GEN_302;
  wire  _GEN_303;
  wire  _GEN_304;
  wire  _GEN_305;
  wire  _GEN_306;
  wire  _GEN_307;
  wire  _GEN_308;
  wire  _GEN_309;
  wire  _GEN_310;
  wire  _GEN_311;
  wire  _GEN_312;
  wire  _GEN_313;
  wire  _GEN_314;
  wire  _GEN_315;
  wire  _GEN_316;
  wire  _GEN_317;
  wire  _GEN_318;
  wire  _GEN_319;
  wire  _GEN_320;
  wire  _GEN_321;
  wire  _GEN_322;
  wire  _GEN_323;
  wire  _GEN_324;
  wire  _GEN_325;
  wire  _GEN_326;
  wire  _GEN_327;
  wire  _GEN_328;
  wire  _GEN_329;
  wire  _GEN_330;
  wire  _GEN_331;
  wire  _GEN_332;
  wire  _GEN_333;
  wire  _GEN_334;
  wire  _GEN_335;
  wire  _GEN_336;
  wire  _GEN_337;
  wire  _GEN_338;
  wire  _GEN_339;
  wire  _GEN_340;
  wire  _GEN_341;
  wire  _GEN_342;
  wire  _GEN_343;
  wire  _GEN_344;
  wire  _GEN_345;
  wire  _GEN_346;
  wire  _GEN_347;
  wire  _GEN_348;
  wire  _GEN_349;
  wire  _GEN_350;
  wire  _GEN_351;
  wire  _GEN_352;
  wire  _GEN_353;
  wire  _GEN_354;
  wire  _GEN_355;
  wire  _GEN_356;
  wire  _GEN_357;
  wire  _GEN_358;
  wire  _GEN_359;
  wire  _GEN_360;
  wire  _GEN_361;
  wire  _GEN_362;
  wire  _GEN_363;
  wire  _GEN_364;
  wire  _GEN_365;
  wire  _GEN_366;
  wire  _GEN_367;
  wire  _GEN_368;
  wire  _GEN_369;
  wire  _GEN_370;
  wire  _GEN_371;
  wire  _GEN_372;
  wire  _GEN_373;
  wire  _GEN_374;
  wire  _GEN_375;
  wire  _GEN_376;
  wire  _GEN_377;
  wire  _GEN_378;
  wire  _GEN_379;
  wire  _GEN_380;
  wire  _GEN_381;
  wire  _GEN_382;
  wire  _GEN_383;
  wire  _GEN_384;
  wire  _GEN_385;
  wire  _GEN_386;
  wire  _GEN_387;
  wire  _GEN_388;
  wire  _GEN_389;
  wire  _GEN_390;
  wire  _GEN_391;
  wire  _GEN_392;
  wire  _GEN_393;
  wire  _GEN_394;
  wire  _GEN_395;
  wire  _GEN_396;
  wire  _GEN_397;
  wire  _GEN_398;
  wire  _GEN_399;
  wire  _GEN_400;
  wire  _GEN_401;
  wire  _GEN_402;
  wire  _GEN_403;
  wire  _GEN_404;
  wire  _GEN_405;
  wire  _GEN_406;
  wire  _GEN_407;
  wire  _GEN_408;
  wire  _GEN_409;
  wire  _GEN_410;
  wire  _GEN_411;
  wire  _GEN_412;
  wire  _GEN_413;
  wire  _GEN_414;
  wire  _GEN_415;
  wire  _GEN_416;
  wire  _GEN_417;
  wire  _GEN_418;
  wire  _GEN_419;
  wire  _GEN_420;
  wire  _GEN_421;
  wire  _GEN_422;
  wire  _GEN_423;
  wire  _GEN_424;
  wire  _GEN_425;
  wire  _GEN_426;
  wire  _GEN_427;
  wire  _GEN_428;
  wire  _GEN_429;
  wire  _GEN_430;
  wire  _GEN_431;
  wire  _GEN_432;
  wire  _GEN_433;
  wire  _GEN_434;
  wire  _GEN_435;
  wire  _GEN_436;
  wire  _GEN_437;
  wire  _GEN_438;
  wire  _GEN_439;
  wire  _GEN_440;
  wire  _GEN_441;
  wire  _GEN_442;
  wire  _GEN_443;
  wire  _GEN_444;
  wire  _GEN_445;
  wire  _GEN_446;
  wire  _GEN_447;
  wire  _GEN_448;
  wire  _GEN_449;
  wire  _GEN_450;
  wire  _GEN_451;
  wire  _GEN_452;
  wire  _GEN_453;
  wire  _GEN_454;
  wire  _GEN_455;
  wire  _GEN_456;
  wire  _GEN_457;
  wire  _GEN_458;
  wire  _GEN_459;
  wire  _GEN_460;
  wire  _GEN_461;
  wire  _GEN_462;
  wire  _GEN_463;
  wire  _GEN_464;
  wire  _GEN_465;
  wire  _GEN_466;
  wire  _GEN_467;
  wire  _GEN_468;
  wire  _GEN_469;
  wire  _GEN_470;
  wire  _GEN_471;
  wire  _GEN_472;
  wire  _GEN_473;
  wire  _GEN_474;
  wire  _GEN_475;
  wire  _GEN_476;
  wire  _GEN_477;
  wire  _GEN_478;
  wire  _GEN_479;
  wire  _GEN_480;
  wire  _GEN_481;
  wire  _GEN_482;
  wire  _GEN_483;
  wire  _GEN_484;
  wire  _GEN_485;
  wire  _GEN_486;
  wire  _GEN_487;
  wire  _GEN_488;
  wire  _GEN_489;
  wire  _GEN_490;
  wire  _GEN_491;
  wire  _GEN_492;
  wire  _GEN_493;
  wire  _GEN_494;
  wire  _GEN_495;
  wire  _GEN_496;
  wire  _GEN_497;
  wire  _GEN_498;
  wire  _GEN_499;
  wire  _GEN_500;
  wire  _GEN_501;
  wire  _GEN_502;
  wire  _GEN_503;
  wire  _GEN_504;
  wire  _GEN_505;
  wire  _GEN_506;
  wire  _GEN_507;
  wire  _GEN_508;
  wire  _GEN_509;
  wire  _GEN_510;
  wire  _GEN_511;
  wire  _GEN_512;
  wire  _T_1053;
  wire  _T_1055;
  wire  _T_1056;
  reg  outputMemBlock_0;
  reg [31:0] _GEN_2052;
  reg  outputMemBlock_1;
  reg [31:0] _GEN_2053;
  reg  outputMemBlock_2;
  reg [31:0] _GEN_2054;
  reg  outputMemBlock_3;
  reg [31:0] _GEN_2055;
  reg  outputMemBlock_4;
  reg [31:0] _GEN_2056;
  reg  outputMemBlock_5;
  reg [31:0] _GEN_2057;
  reg  outputMemBlock_6;
  reg [31:0] _GEN_2058;
  reg  outputMemBlock_7;
  reg [31:0] _GEN_2059;
  reg  outputMemBlock_8;
  reg [31:0] _GEN_2060;
  reg  outputMemBlock_9;
  reg [31:0] _GEN_2061;
  reg  outputMemBlock_10;
  reg [31:0] _GEN_2062;
  reg  outputMemBlock_11;
  reg [31:0] _GEN_2063;
  reg  outputMemBlock_12;
  reg [31:0] _GEN_2064;
  reg  outputMemBlock_13;
  reg [31:0] _GEN_2065;
  reg  outputMemBlock_14;
  reg [31:0] _GEN_2066;
  reg  outputMemBlock_15;
  reg [31:0] _GEN_2067;
  reg  outputMemBlock_16;
  reg [31:0] _GEN_2068;
  reg  outputMemBlock_17;
  reg [31:0] _GEN_2069;
  reg  outputMemBlock_18;
  reg [31:0] _GEN_2070;
  reg  outputMemBlock_19;
  reg [31:0] _GEN_2071;
  reg  outputMemBlock_20;
  reg [31:0] _GEN_2072;
  reg  outputMemBlock_21;
  reg [31:0] _GEN_2073;
  reg  outputMemBlock_22;
  reg [31:0] _GEN_2074;
  reg  outputMemBlock_23;
  reg [31:0] _GEN_2075;
  reg  outputMemBlock_24;
  reg [31:0] _GEN_2076;
  reg  outputMemBlock_25;
  reg [31:0] _GEN_2077;
  reg  outputMemBlock_26;
  reg [31:0] _GEN_2078;
  reg  outputMemBlock_27;
  reg [31:0] _GEN_2079;
  reg  outputMemBlock_28;
  reg [31:0] _GEN_2080;
  reg  outputMemBlock_29;
  reg [31:0] _GEN_2081;
  reg  outputMemBlock_30;
  reg [31:0] _GEN_2082;
  reg  outputMemBlock_31;
  reg [31:0] _GEN_2083;
  reg  outputMemBlock_32;
  reg [31:0] _GEN_2084;
  reg  outputMemBlock_33;
  reg [31:0] _GEN_2085;
  reg  outputMemBlock_34;
  reg [31:0] _GEN_2086;
  reg  outputMemBlock_35;
  reg [31:0] _GEN_2087;
  reg  outputMemBlock_36;
  reg [31:0] _GEN_2088;
  reg  outputMemBlock_37;
  reg [31:0] _GEN_2089;
  reg  outputMemBlock_38;
  reg [31:0] _GEN_2090;
  reg  outputMemBlock_39;
  reg [31:0] _GEN_2091;
  reg  outputMemBlock_40;
  reg [31:0] _GEN_2092;
  reg  outputMemBlock_41;
  reg [31:0] _GEN_2093;
  reg  outputMemBlock_42;
  reg [31:0] _GEN_2094;
  reg  outputMemBlock_43;
  reg [31:0] _GEN_2095;
  reg  outputMemBlock_44;
  reg [31:0] _GEN_2096;
  reg  outputMemBlock_45;
  reg [31:0] _GEN_2097;
  reg  outputMemBlock_46;
  reg [31:0] _GEN_2098;
  reg  outputMemBlock_47;
  reg [31:0] _GEN_2099;
  reg  outputMemBlock_48;
  reg [31:0] _GEN_2100;
  reg  outputMemBlock_49;
  reg [31:0] _GEN_2101;
  reg  outputMemBlock_50;
  reg [31:0] _GEN_2102;
  reg  outputMemBlock_51;
  reg [31:0] _GEN_2103;
  reg  outputMemBlock_52;
  reg [31:0] _GEN_2104;
  reg  outputMemBlock_53;
  reg [31:0] _GEN_2105;
  reg  outputMemBlock_54;
  reg [31:0] _GEN_2106;
  reg  outputMemBlock_55;
  reg [31:0] _GEN_2107;
  reg  outputMemBlock_56;
  reg [31:0] _GEN_2108;
  reg  outputMemBlock_57;
  reg [31:0] _GEN_2109;
  reg  outputMemBlock_58;
  reg [31:0] _GEN_2110;
  reg  outputMemBlock_59;
  reg [31:0] _GEN_2111;
  reg  outputMemBlock_60;
  reg [31:0] _GEN_2112;
  reg  outputMemBlock_61;
  reg [31:0] _GEN_2113;
  reg  outputMemBlock_62;
  reg [31:0] _GEN_2114;
  reg  outputMemBlock_63;
  reg [31:0] _GEN_2115;
  reg  outputMemBlock_64;
  reg [31:0] _GEN_2116;
  reg  outputMemBlock_65;
  reg [31:0] _GEN_2117;
  reg  outputMemBlock_66;
  reg [31:0] _GEN_2118;
  reg  outputMemBlock_67;
  reg [31:0] _GEN_2119;
  reg  outputMemBlock_68;
  reg [31:0] _GEN_2120;
  reg  outputMemBlock_69;
  reg [31:0] _GEN_2121;
  reg  outputMemBlock_70;
  reg [31:0] _GEN_2122;
  reg  outputMemBlock_71;
  reg [31:0] _GEN_2123;
  reg  outputMemBlock_72;
  reg [31:0] _GEN_2124;
  reg  outputMemBlock_73;
  reg [31:0] _GEN_2125;
  reg  outputMemBlock_74;
  reg [31:0] _GEN_2126;
  reg  outputMemBlock_75;
  reg [31:0] _GEN_2127;
  reg  outputMemBlock_76;
  reg [31:0] _GEN_2128;
  reg  outputMemBlock_77;
  reg [31:0] _GEN_2129;
  reg  outputMemBlock_78;
  reg [31:0] _GEN_2130;
  reg  outputMemBlock_79;
  reg [31:0] _GEN_2131;
  reg  outputMemBlock_80;
  reg [31:0] _GEN_2132;
  reg  outputMemBlock_81;
  reg [31:0] _GEN_2133;
  reg  outputMemBlock_82;
  reg [31:0] _GEN_2134;
  reg  outputMemBlock_83;
  reg [31:0] _GEN_2135;
  reg  outputMemBlock_84;
  reg [31:0] _GEN_2136;
  reg  outputMemBlock_85;
  reg [31:0] _GEN_2137;
  reg  outputMemBlock_86;
  reg [31:0] _GEN_2138;
  reg  outputMemBlock_87;
  reg [31:0] _GEN_2139;
  reg  outputMemBlock_88;
  reg [31:0] _GEN_2140;
  reg  outputMemBlock_89;
  reg [31:0] _GEN_2141;
  reg  outputMemBlock_90;
  reg [31:0] _GEN_2142;
  reg  outputMemBlock_91;
  reg [31:0] _GEN_2143;
  reg  outputMemBlock_92;
  reg [31:0] _GEN_2144;
  reg  outputMemBlock_93;
  reg [31:0] _GEN_2145;
  reg  outputMemBlock_94;
  reg [31:0] _GEN_2146;
  reg  outputMemBlock_95;
  reg [31:0] _GEN_2147;
  reg  outputMemBlock_96;
  reg [31:0] _GEN_2148;
  reg  outputMemBlock_97;
  reg [31:0] _GEN_2149;
  reg  outputMemBlock_98;
  reg [31:0] _GEN_2150;
  reg  outputMemBlock_99;
  reg [31:0] _GEN_2151;
  reg  outputMemBlock_100;
  reg [31:0] _GEN_2152;
  reg  outputMemBlock_101;
  reg [31:0] _GEN_2153;
  reg  outputMemBlock_102;
  reg [31:0] _GEN_2154;
  reg  outputMemBlock_103;
  reg [31:0] _GEN_2155;
  reg  outputMemBlock_104;
  reg [31:0] _GEN_2156;
  reg  outputMemBlock_105;
  reg [31:0] _GEN_2157;
  reg  outputMemBlock_106;
  reg [31:0] _GEN_2158;
  reg  outputMemBlock_107;
  reg [31:0] _GEN_2159;
  reg  outputMemBlock_108;
  reg [31:0] _GEN_2160;
  reg  outputMemBlock_109;
  reg [31:0] _GEN_2161;
  reg  outputMemBlock_110;
  reg [31:0] _GEN_2162;
  reg  outputMemBlock_111;
  reg [31:0] _GEN_2163;
  reg  outputMemBlock_112;
  reg [31:0] _GEN_2164;
  reg  outputMemBlock_113;
  reg [31:0] _GEN_2165;
  reg  outputMemBlock_114;
  reg [31:0] _GEN_2166;
  reg  outputMemBlock_115;
  reg [31:0] _GEN_2167;
  reg  outputMemBlock_116;
  reg [31:0] _GEN_2168;
  reg  outputMemBlock_117;
  reg [31:0] _GEN_2169;
  reg  outputMemBlock_118;
  reg [31:0] _GEN_2170;
  reg  outputMemBlock_119;
  reg [31:0] _GEN_2171;
  reg  outputMemBlock_120;
  reg [31:0] _GEN_2172;
  reg  outputMemBlock_121;
  reg [31:0] _GEN_2173;
  reg  outputMemBlock_122;
  reg [31:0] _GEN_2174;
  reg  outputMemBlock_123;
  reg [31:0] _GEN_2175;
  reg  outputMemBlock_124;
  reg [31:0] _GEN_2176;
  reg  outputMemBlock_125;
  reg [31:0] _GEN_2177;
  reg  outputMemBlock_126;
  reg [31:0] _GEN_2178;
  reg  outputMemBlock_127;
  reg [31:0] _GEN_2179;
  reg  outputMemBlock_128;
  reg [31:0] _GEN_2180;
  reg  outputMemBlock_129;
  reg [31:0] _GEN_2181;
  reg  outputMemBlock_130;
  reg [31:0] _GEN_2182;
  reg  outputMemBlock_131;
  reg [31:0] _GEN_2183;
  reg  outputMemBlock_132;
  reg [31:0] _GEN_2184;
  reg  outputMemBlock_133;
  reg [31:0] _GEN_2185;
  reg  outputMemBlock_134;
  reg [31:0] _GEN_2186;
  reg  outputMemBlock_135;
  reg [31:0] _GEN_2187;
  reg  outputMemBlock_136;
  reg [31:0] _GEN_2188;
  reg  outputMemBlock_137;
  reg [31:0] _GEN_2189;
  reg  outputMemBlock_138;
  reg [31:0] _GEN_2190;
  reg  outputMemBlock_139;
  reg [31:0] _GEN_2191;
  reg  outputMemBlock_140;
  reg [31:0] _GEN_2192;
  reg  outputMemBlock_141;
  reg [31:0] _GEN_2193;
  reg  outputMemBlock_142;
  reg [31:0] _GEN_2194;
  reg  outputMemBlock_143;
  reg [31:0] _GEN_2195;
  reg  outputMemBlock_144;
  reg [31:0] _GEN_2196;
  reg  outputMemBlock_145;
  reg [31:0] _GEN_2197;
  reg  outputMemBlock_146;
  reg [31:0] _GEN_2198;
  reg  outputMemBlock_147;
  reg [31:0] _GEN_2199;
  reg  outputMemBlock_148;
  reg [31:0] _GEN_2200;
  reg  outputMemBlock_149;
  reg [31:0] _GEN_2201;
  reg  outputMemBlock_150;
  reg [31:0] _GEN_2202;
  reg  outputMemBlock_151;
  reg [31:0] _GEN_2203;
  reg  outputMemBlock_152;
  reg [31:0] _GEN_2204;
  reg  outputMemBlock_153;
  reg [31:0] _GEN_2205;
  reg  outputMemBlock_154;
  reg [31:0] _GEN_2206;
  reg  outputMemBlock_155;
  reg [31:0] _GEN_2207;
  reg  outputMemBlock_156;
  reg [31:0] _GEN_2208;
  reg  outputMemBlock_157;
  reg [31:0] _GEN_2209;
  reg  outputMemBlock_158;
  reg [31:0] _GEN_2210;
  reg  outputMemBlock_159;
  reg [31:0] _GEN_2211;
  reg  outputMemBlock_160;
  reg [31:0] _GEN_2212;
  reg  outputMemBlock_161;
  reg [31:0] _GEN_2213;
  reg  outputMemBlock_162;
  reg [31:0] _GEN_2214;
  reg  outputMemBlock_163;
  reg [31:0] _GEN_2215;
  reg  outputMemBlock_164;
  reg [31:0] _GEN_2216;
  reg  outputMemBlock_165;
  reg [31:0] _GEN_2217;
  reg  outputMemBlock_166;
  reg [31:0] _GEN_2218;
  reg  outputMemBlock_167;
  reg [31:0] _GEN_2219;
  reg  outputMemBlock_168;
  reg [31:0] _GEN_2220;
  reg  outputMemBlock_169;
  reg [31:0] _GEN_2221;
  reg  outputMemBlock_170;
  reg [31:0] _GEN_2222;
  reg  outputMemBlock_171;
  reg [31:0] _GEN_2223;
  reg  outputMemBlock_172;
  reg [31:0] _GEN_2224;
  reg  outputMemBlock_173;
  reg [31:0] _GEN_2225;
  reg  outputMemBlock_174;
  reg [31:0] _GEN_2226;
  reg  outputMemBlock_175;
  reg [31:0] _GEN_2227;
  reg  outputMemBlock_176;
  reg [31:0] _GEN_2228;
  reg  outputMemBlock_177;
  reg [31:0] _GEN_2229;
  reg  outputMemBlock_178;
  reg [31:0] _GEN_2230;
  reg  outputMemBlock_179;
  reg [31:0] _GEN_2231;
  reg  outputMemBlock_180;
  reg [31:0] _GEN_2232;
  reg  outputMemBlock_181;
  reg [31:0] _GEN_2233;
  reg  outputMemBlock_182;
  reg [31:0] _GEN_2234;
  reg  outputMemBlock_183;
  reg [31:0] _GEN_2235;
  reg  outputMemBlock_184;
  reg [31:0] _GEN_2236;
  reg  outputMemBlock_185;
  reg [31:0] _GEN_2237;
  reg  outputMemBlock_186;
  reg [31:0] _GEN_2238;
  reg  outputMemBlock_187;
  reg [31:0] _GEN_2239;
  reg  outputMemBlock_188;
  reg [31:0] _GEN_2240;
  reg  outputMemBlock_189;
  reg [31:0] _GEN_2241;
  reg  outputMemBlock_190;
  reg [31:0] _GEN_2242;
  reg  outputMemBlock_191;
  reg [31:0] _GEN_2243;
  reg  outputMemBlock_192;
  reg [31:0] _GEN_2244;
  reg  outputMemBlock_193;
  reg [31:0] _GEN_2245;
  reg  outputMemBlock_194;
  reg [31:0] _GEN_2246;
  reg  outputMemBlock_195;
  reg [31:0] _GEN_2247;
  reg  outputMemBlock_196;
  reg [31:0] _GEN_2248;
  reg  outputMemBlock_197;
  reg [31:0] _GEN_2249;
  reg  outputMemBlock_198;
  reg [31:0] _GEN_2250;
  reg  outputMemBlock_199;
  reg [31:0] _GEN_2251;
  reg  outputMemBlock_200;
  reg [31:0] _GEN_2252;
  reg  outputMemBlock_201;
  reg [31:0] _GEN_2253;
  reg  outputMemBlock_202;
  reg [31:0] _GEN_2254;
  reg  outputMemBlock_203;
  reg [31:0] _GEN_2255;
  reg  outputMemBlock_204;
  reg [31:0] _GEN_2256;
  reg  outputMemBlock_205;
  reg [31:0] _GEN_2257;
  reg  outputMemBlock_206;
  reg [31:0] _GEN_2258;
  reg  outputMemBlock_207;
  reg [31:0] _GEN_2259;
  reg  outputMemBlock_208;
  reg [31:0] _GEN_2260;
  reg  outputMemBlock_209;
  reg [31:0] _GEN_2261;
  reg  outputMemBlock_210;
  reg [31:0] _GEN_2262;
  reg  outputMemBlock_211;
  reg [31:0] _GEN_2263;
  reg  outputMemBlock_212;
  reg [31:0] _GEN_2264;
  reg  outputMemBlock_213;
  reg [31:0] _GEN_2265;
  reg  outputMemBlock_214;
  reg [31:0] _GEN_2266;
  reg  outputMemBlock_215;
  reg [31:0] _GEN_2267;
  reg  outputMemBlock_216;
  reg [31:0] _GEN_2268;
  reg  outputMemBlock_217;
  reg [31:0] _GEN_2269;
  reg  outputMemBlock_218;
  reg [31:0] _GEN_2270;
  reg  outputMemBlock_219;
  reg [31:0] _GEN_2271;
  reg  outputMemBlock_220;
  reg [31:0] _GEN_2272;
  reg  outputMemBlock_221;
  reg [31:0] _GEN_2273;
  reg  outputMemBlock_222;
  reg [31:0] _GEN_2274;
  reg  outputMemBlock_223;
  reg [31:0] _GEN_2275;
  reg  outputMemBlock_224;
  reg [31:0] _GEN_2276;
  reg  outputMemBlock_225;
  reg [31:0] _GEN_2277;
  reg  outputMemBlock_226;
  reg [31:0] _GEN_2278;
  reg  outputMemBlock_227;
  reg [31:0] _GEN_2279;
  reg  outputMemBlock_228;
  reg [31:0] _GEN_2280;
  reg  outputMemBlock_229;
  reg [31:0] _GEN_2281;
  reg  outputMemBlock_230;
  reg [31:0] _GEN_2282;
  reg  outputMemBlock_231;
  reg [31:0] _GEN_2283;
  reg  outputMemBlock_232;
  reg [31:0] _GEN_2284;
  reg  outputMemBlock_233;
  reg [31:0] _GEN_2285;
  reg  outputMemBlock_234;
  reg [31:0] _GEN_2286;
  reg  outputMemBlock_235;
  reg [31:0] _GEN_2287;
  reg  outputMemBlock_236;
  reg [31:0] _GEN_2288;
  reg  outputMemBlock_237;
  reg [31:0] _GEN_2289;
  reg  outputMemBlock_238;
  reg [31:0] _GEN_2290;
  reg  outputMemBlock_239;
  reg [31:0] _GEN_2291;
  reg  outputMemBlock_240;
  reg [31:0] _GEN_2292;
  reg  outputMemBlock_241;
  reg [31:0] _GEN_2293;
  reg  outputMemBlock_242;
  reg [31:0] _GEN_2294;
  reg  outputMemBlock_243;
  reg [31:0] _GEN_2295;
  reg  outputMemBlock_244;
  reg [31:0] _GEN_2296;
  reg  outputMemBlock_245;
  reg [31:0] _GEN_2297;
  reg  outputMemBlock_246;
  reg [31:0] _GEN_2298;
  reg  outputMemBlock_247;
  reg [31:0] _GEN_2299;
  reg  outputMemBlock_248;
  reg [31:0] _GEN_2300;
  reg  outputMemBlock_249;
  reg [31:0] _GEN_2301;
  reg  outputMemBlock_250;
  reg [31:0] _GEN_2302;
  reg  outputMemBlock_251;
  reg [31:0] _GEN_2303;
  reg  outputMemBlock_252;
  reg [31:0] _GEN_2304;
  reg  outputMemBlock_253;
  reg [31:0] _GEN_2305;
  reg  outputMemBlock_254;
  reg [31:0] _GEN_2306;
  reg  outputMemBlock_255;
  reg [31:0] _GEN_2307;
  reg  outputMemBlock_256;
  reg [31:0] _GEN_2308;
  reg  outputMemBlock_257;
  reg [31:0] _GEN_2309;
  reg  outputMemBlock_258;
  reg [31:0] _GEN_2310;
  reg  outputMemBlock_259;
  reg [31:0] _GEN_2311;
  reg  outputMemBlock_260;
  reg [31:0] _GEN_2312;
  reg  outputMemBlock_261;
  reg [31:0] _GEN_2313;
  reg  outputMemBlock_262;
  reg [31:0] _GEN_2314;
  reg  outputMemBlock_263;
  reg [31:0] _GEN_2315;
  reg  outputMemBlock_264;
  reg [31:0] _GEN_2316;
  reg  outputMemBlock_265;
  reg [31:0] _GEN_2317;
  reg  outputMemBlock_266;
  reg [31:0] _GEN_2318;
  reg  outputMemBlock_267;
  reg [31:0] _GEN_2319;
  reg  outputMemBlock_268;
  reg [31:0] _GEN_2320;
  reg  outputMemBlock_269;
  reg [31:0] _GEN_2321;
  reg  outputMemBlock_270;
  reg [31:0] _GEN_2322;
  reg  outputMemBlock_271;
  reg [31:0] _GEN_2323;
  reg  outputMemBlock_272;
  reg [31:0] _GEN_2324;
  reg  outputMemBlock_273;
  reg [31:0] _GEN_2325;
  reg  outputMemBlock_274;
  reg [31:0] _GEN_2326;
  reg  outputMemBlock_275;
  reg [31:0] _GEN_2327;
  reg  outputMemBlock_276;
  reg [31:0] _GEN_2328;
  reg  outputMemBlock_277;
  reg [31:0] _GEN_2329;
  reg  outputMemBlock_278;
  reg [31:0] _GEN_2330;
  reg  outputMemBlock_279;
  reg [31:0] _GEN_2331;
  reg  outputMemBlock_280;
  reg [31:0] _GEN_2332;
  reg  outputMemBlock_281;
  reg [31:0] _GEN_2333;
  reg  outputMemBlock_282;
  reg [31:0] _GEN_2334;
  reg  outputMemBlock_283;
  reg [31:0] _GEN_2335;
  reg  outputMemBlock_284;
  reg [31:0] _GEN_2336;
  reg  outputMemBlock_285;
  reg [31:0] _GEN_2337;
  reg  outputMemBlock_286;
  reg [31:0] _GEN_2338;
  reg  outputMemBlock_287;
  reg [31:0] _GEN_2339;
  reg  outputMemBlock_288;
  reg [31:0] _GEN_2340;
  reg  outputMemBlock_289;
  reg [31:0] _GEN_2341;
  reg  outputMemBlock_290;
  reg [31:0] _GEN_2342;
  reg  outputMemBlock_291;
  reg [31:0] _GEN_2343;
  reg  outputMemBlock_292;
  reg [31:0] _GEN_2344;
  reg  outputMemBlock_293;
  reg [31:0] _GEN_2345;
  reg  outputMemBlock_294;
  reg [31:0] _GEN_2346;
  reg  outputMemBlock_295;
  reg [31:0] _GEN_2347;
  reg  outputMemBlock_296;
  reg [31:0] _GEN_2348;
  reg  outputMemBlock_297;
  reg [31:0] _GEN_2349;
  reg  outputMemBlock_298;
  reg [31:0] _GEN_2350;
  reg  outputMemBlock_299;
  reg [31:0] _GEN_2351;
  reg  outputMemBlock_300;
  reg [31:0] _GEN_2352;
  reg  outputMemBlock_301;
  reg [31:0] _GEN_2353;
  reg  outputMemBlock_302;
  reg [31:0] _GEN_2354;
  reg  outputMemBlock_303;
  reg [31:0] _GEN_2355;
  reg  outputMemBlock_304;
  reg [31:0] _GEN_2356;
  reg  outputMemBlock_305;
  reg [31:0] _GEN_2357;
  reg  outputMemBlock_306;
  reg [31:0] _GEN_2358;
  reg  outputMemBlock_307;
  reg [31:0] _GEN_2359;
  reg  outputMemBlock_308;
  reg [31:0] _GEN_2360;
  reg  outputMemBlock_309;
  reg [31:0] _GEN_2361;
  reg  outputMemBlock_310;
  reg [31:0] _GEN_2362;
  reg  outputMemBlock_311;
  reg [31:0] _GEN_2363;
  reg  outputMemBlock_312;
  reg [31:0] _GEN_2364;
  reg  outputMemBlock_313;
  reg [31:0] _GEN_2365;
  reg  outputMemBlock_314;
  reg [31:0] _GEN_2366;
  reg  outputMemBlock_315;
  reg [31:0] _GEN_2367;
  reg  outputMemBlock_316;
  reg [31:0] _GEN_2368;
  reg  outputMemBlock_317;
  reg [31:0] _GEN_2369;
  reg  outputMemBlock_318;
  reg [31:0] _GEN_2370;
  reg  outputMemBlock_319;
  reg [31:0] _GEN_2371;
  reg  outputMemBlock_320;
  reg [31:0] _GEN_2372;
  reg  outputMemBlock_321;
  reg [31:0] _GEN_2373;
  reg  outputMemBlock_322;
  reg [31:0] _GEN_2374;
  reg  outputMemBlock_323;
  reg [31:0] _GEN_2375;
  reg  outputMemBlock_324;
  reg [31:0] _GEN_2376;
  reg  outputMemBlock_325;
  reg [31:0] _GEN_2377;
  reg  outputMemBlock_326;
  reg [31:0] _GEN_2378;
  reg  outputMemBlock_327;
  reg [31:0] _GEN_2379;
  reg  outputMemBlock_328;
  reg [31:0] _GEN_2380;
  reg  outputMemBlock_329;
  reg [31:0] _GEN_2381;
  reg  outputMemBlock_330;
  reg [31:0] _GEN_2382;
  reg  outputMemBlock_331;
  reg [31:0] _GEN_2383;
  reg  outputMemBlock_332;
  reg [31:0] _GEN_2384;
  reg  outputMemBlock_333;
  reg [31:0] _GEN_2385;
  reg  outputMemBlock_334;
  reg [31:0] _GEN_2386;
  reg  outputMemBlock_335;
  reg [31:0] _GEN_2387;
  reg  outputMemBlock_336;
  reg [31:0] _GEN_2388;
  reg  outputMemBlock_337;
  reg [31:0] _GEN_2389;
  reg  outputMemBlock_338;
  reg [31:0] _GEN_2390;
  reg  outputMemBlock_339;
  reg [31:0] _GEN_2391;
  reg  outputMemBlock_340;
  reg [31:0] _GEN_2392;
  reg  outputMemBlock_341;
  reg [31:0] _GEN_2393;
  reg  outputMemBlock_342;
  reg [31:0] _GEN_2394;
  reg  outputMemBlock_343;
  reg [31:0] _GEN_2395;
  reg  outputMemBlock_344;
  reg [31:0] _GEN_2396;
  reg  outputMemBlock_345;
  reg [31:0] _GEN_2397;
  reg  outputMemBlock_346;
  reg [31:0] _GEN_2398;
  reg  outputMemBlock_347;
  reg [31:0] _GEN_2399;
  reg  outputMemBlock_348;
  reg [31:0] _GEN_2400;
  reg  outputMemBlock_349;
  reg [31:0] _GEN_2401;
  reg  outputMemBlock_350;
  reg [31:0] _GEN_2402;
  reg  outputMemBlock_351;
  reg [31:0] _GEN_2403;
  reg  outputMemBlock_352;
  reg [31:0] _GEN_2404;
  reg  outputMemBlock_353;
  reg [31:0] _GEN_2405;
  reg  outputMemBlock_354;
  reg [31:0] _GEN_2406;
  reg  outputMemBlock_355;
  reg [31:0] _GEN_2407;
  reg  outputMemBlock_356;
  reg [31:0] _GEN_2408;
  reg  outputMemBlock_357;
  reg [31:0] _GEN_2409;
  reg  outputMemBlock_358;
  reg [31:0] _GEN_2410;
  reg  outputMemBlock_359;
  reg [31:0] _GEN_2411;
  reg  outputMemBlock_360;
  reg [31:0] _GEN_2412;
  reg  outputMemBlock_361;
  reg [31:0] _GEN_2413;
  reg  outputMemBlock_362;
  reg [31:0] _GEN_2414;
  reg  outputMemBlock_363;
  reg [31:0] _GEN_2415;
  reg  outputMemBlock_364;
  reg [31:0] _GEN_2416;
  reg  outputMemBlock_365;
  reg [31:0] _GEN_2417;
  reg  outputMemBlock_366;
  reg [31:0] _GEN_2418;
  reg  outputMemBlock_367;
  reg [31:0] _GEN_2419;
  reg  outputMemBlock_368;
  reg [31:0] _GEN_2420;
  reg  outputMemBlock_369;
  reg [31:0] _GEN_2421;
  reg  outputMemBlock_370;
  reg [31:0] _GEN_2422;
  reg  outputMemBlock_371;
  reg [31:0] _GEN_2423;
  reg  outputMemBlock_372;
  reg [31:0] _GEN_2424;
  reg  outputMemBlock_373;
  reg [31:0] _GEN_2425;
  reg  outputMemBlock_374;
  reg [31:0] _GEN_2426;
  reg  outputMemBlock_375;
  reg [31:0] _GEN_2427;
  reg  outputMemBlock_376;
  reg [31:0] _GEN_2428;
  reg  outputMemBlock_377;
  reg [31:0] _GEN_2429;
  reg  outputMemBlock_378;
  reg [31:0] _GEN_2430;
  reg  outputMemBlock_379;
  reg [31:0] _GEN_2431;
  reg  outputMemBlock_380;
  reg [31:0] _GEN_2432;
  reg  outputMemBlock_381;
  reg [31:0] _GEN_2433;
  reg  outputMemBlock_382;
  reg [31:0] _GEN_2434;
  reg  outputMemBlock_383;
  reg [31:0] _GEN_2435;
  reg  outputMemBlock_384;
  reg [31:0] _GEN_2436;
  reg  outputMemBlock_385;
  reg [31:0] _GEN_2437;
  reg  outputMemBlock_386;
  reg [31:0] _GEN_2438;
  reg  outputMemBlock_387;
  reg [31:0] _GEN_2439;
  reg  outputMemBlock_388;
  reg [31:0] _GEN_2440;
  reg  outputMemBlock_389;
  reg [31:0] _GEN_2441;
  reg  outputMemBlock_390;
  reg [31:0] _GEN_2442;
  reg  outputMemBlock_391;
  reg [31:0] _GEN_2443;
  reg  outputMemBlock_392;
  reg [31:0] _GEN_2444;
  reg  outputMemBlock_393;
  reg [31:0] _GEN_2445;
  reg  outputMemBlock_394;
  reg [31:0] _GEN_2446;
  reg  outputMemBlock_395;
  reg [31:0] _GEN_2447;
  reg  outputMemBlock_396;
  reg [31:0] _GEN_2448;
  reg  outputMemBlock_397;
  reg [31:0] _GEN_2449;
  reg  outputMemBlock_398;
  reg [31:0] _GEN_2450;
  reg  outputMemBlock_399;
  reg [31:0] _GEN_2451;
  reg  outputMemBlock_400;
  reg [31:0] _GEN_2452;
  reg  outputMemBlock_401;
  reg [31:0] _GEN_2453;
  reg  outputMemBlock_402;
  reg [31:0] _GEN_2454;
  reg  outputMemBlock_403;
  reg [31:0] _GEN_2455;
  reg  outputMemBlock_404;
  reg [31:0] _GEN_2456;
  reg  outputMemBlock_405;
  reg [31:0] _GEN_2457;
  reg  outputMemBlock_406;
  reg [31:0] _GEN_2458;
  reg  outputMemBlock_407;
  reg [31:0] _GEN_2459;
  reg  outputMemBlock_408;
  reg [31:0] _GEN_2460;
  reg  outputMemBlock_409;
  reg [31:0] _GEN_2461;
  reg  outputMemBlock_410;
  reg [31:0] _GEN_2462;
  reg  outputMemBlock_411;
  reg [31:0] _GEN_2463;
  reg  outputMemBlock_412;
  reg [31:0] _GEN_2464;
  reg  outputMemBlock_413;
  reg [31:0] _GEN_2465;
  reg  outputMemBlock_414;
  reg [31:0] _GEN_2466;
  reg  outputMemBlock_415;
  reg [31:0] _GEN_2467;
  reg  outputMemBlock_416;
  reg [31:0] _GEN_2468;
  reg  outputMemBlock_417;
  reg [31:0] _GEN_2469;
  reg  outputMemBlock_418;
  reg [31:0] _GEN_2470;
  reg  outputMemBlock_419;
  reg [31:0] _GEN_2471;
  reg  outputMemBlock_420;
  reg [31:0] _GEN_2472;
  reg  outputMemBlock_421;
  reg [31:0] _GEN_2473;
  reg  outputMemBlock_422;
  reg [31:0] _GEN_2474;
  reg  outputMemBlock_423;
  reg [31:0] _GEN_2475;
  reg  outputMemBlock_424;
  reg [31:0] _GEN_2476;
  reg  outputMemBlock_425;
  reg [31:0] _GEN_2477;
  reg  outputMemBlock_426;
  reg [31:0] _GEN_2478;
  reg  outputMemBlock_427;
  reg [31:0] _GEN_2479;
  reg  outputMemBlock_428;
  reg [31:0] _GEN_2480;
  reg  outputMemBlock_429;
  reg [31:0] _GEN_2481;
  reg  outputMemBlock_430;
  reg [31:0] _GEN_2482;
  reg  outputMemBlock_431;
  reg [31:0] _GEN_2483;
  reg  outputMemBlock_432;
  reg [31:0] _GEN_2484;
  reg  outputMemBlock_433;
  reg [31:0] _GEN_2485;
  reg  outputMemBlock_434;
  reg [31:0] _GEN_2486;
  reg  outputMemBlock_435;
  reg [31:0] _GEN_2487;
  reg  outputMemBlock_436;
  reg [31:0] _GEN_2488;
  reg  outputMemBlock_437;
  reg [31:0] _GEN_2489;
  reg  outputMemBlock_438;
  reg [31:0] _GEN_2490;
  reg  outputMemBlock_439;
  reg [31:0] _GEN_2491;
  reg  outputMemBlock_440;
  reg [31:0] _GEN_2492;
  reg  outputMemBlock_441;
  reg [31:0] _GEN_2493;
  reg  outputMemBlock_442;
  reg [31:0] _GEN_2494;
  reg  outputMemBlock_443;
  reg [31:0] _GEN_2495;
  reg  outputMemBlock_444;
  reg [31:0] _GEN_2496;
  reg  outputMemBlock_445;
  reg [31:0] _GEN_2497;
  reg  outputMemBlock_446;
  reg [31:0] _GEN_2498;
  reg  outputMemBlock_447;
  reg [31:0] _GEN_2499;
  reg  outputMemBlock_448;
  reg [31:0] _GEN_2500;
  reg  outputMemBlock_449;
  reg [31:0] _GEN_2501;
  reg  outputMemBlock_450;
  reg [31:0] _GEN_2502;
  reg  outputMemBlock_451;
  reg [31:0] _GEN_2503;
  reg  outputMemBlock_452;
  reg [31:0] _GEN_2504;
  reg  outputMemBlock_453;
  reg [31:0] _GEN_2505;
  reg  outputMemBlock_454;
  reg [31:0] _GEN_2506;
  reg  outputMemBlock_455;
  reg [31:0] _GEN_2507;
  reg  outputMemBlock_456;
  reg [31:0] _GEN_2508;
  reg  outputMemBlock_457;
  reg [31:0] _GEN_2509;
  reg  outputMemBlock_458;
  reg [31:0] _GEN_2510;
  reg  outputMemBlock_459;
  reg [31:0] _GEN_2511;
  reg  outputMemBlock_460;
  reg [31:0] _GEN_2512;
  reg  outputMemBlock_461;
  reg [31:0] _GEN_2513;
  reg  outputMemBlock_462;
  reg [31:0] _GEN_2514;
  reg  outputMemBlock_463;
  reg [31:0] _GEN_2515;
  reg  outputMemBlock_464;
  reg [31:0] _GEN_2516;
  reg  outputMemBlock_465;
  reg [31:0] _GEN_2517;
  reg  outputMemBlock_466;
  reg [31:0] _GEN_2518;
  reg  outputMemBlock_467;
  reg [31:0] _GEN_2519;
  reg  outputMemBlock_468;
  reg [31:0] _GEN_2520;
  reg  outputMemBlock_469;
  reg [31:0] _GEN_2521;
  reg  outputMemBlock_470;
  reg [31:0] _GEN_2522;
  reg  outputMemBlock_471;
  reg [31:0] _GEN_2523;
  reg  outputMemBlock_472;
  reg [31:0] _GEN_2524;
  reg  outputMemBlock_473;
  reg [31:0] _GEN_2525;
  reg  outputMemBlock_474;
  reg [31:0] _GEN_2526;
  reg  outputMemBlock_475;
  reg [31:0] _GEN_2527;
  reg  outputMemBlock_476;
  reg [31:0] _GEN_2528;
  reg  outputMemBlock_477;
  reg [31:0] _GEN_2529;
  reg  outputMemBlock_478;
  reg [31:0] _GEN_2530;
  reg  outputMemBlock_479;
  reg [31:0] _GEN_2531;
  reg  outputMemBlock_480;
  reg [31:0] _GEN_2532;
  reg  outputMemBlock_481;
  reg [31:0] _GEN_2533;
  reg  outputMemBlock_482;
  reg [31:0] _GEN_2534;
  reg  outputMemBlock_483;
  reg [31:0] _GEN_2535;
  reg  outputMemBlock_484;
  reg [31:0] _GEN_2536;
  reg  outputMemBlock_485;
  reg [31:0] _GEN_2537;
  reg  outputMemBlock_486;
  reg [31:0] _GEN_2538;
  reg  outputMemBlock_487;
  reg [31:0] _GEN_2539;
  reg  outputMemBlock_488;
  reg [31:0] _GEN_2540;
  reg  outputMemBlock_489;
  reg [31:0] _GEN_2541;
  reg  outputMemBlock_490;
  reg [31:0] _GEN_2542;
  reg  outputMemBlock_491;
  reg [31:0] _GEN_2543;
  reg  outputMemBlock_492;
  reg [31:0] _GEN_2544;
  reg  outputMemBlock_493;
  reg [31:0] _GEN_2545;
  reg  outputMemBlock_494;
  reg [31:0] _GEN_2546;
  reg  outputMemBlock_495;
  reg [31:0] _GEN_2547;
  reg  outputMemBlock_496;
  reg [31:0] _GEN_2548;
  reg  outputMemBlock_497;
  reg [31:0] _GEN_2549;
  reg  outputMemBlock_498;
  reg [31:0] _GEN_2550;
  reg  outputMemBlock_499;
  reg [31:0] _GEN_2551;
  reg  outputMemBlock_500;
  reg [31:0] _GEN_2552;
  reg  outputMemBlock_501;
  reg [31:0] _GEN_2553;
  reg  outputMemBlock_502;
  reg [31:0] _GEN_2554;
  reg  outputMemBlock_503;
  reg [31:0] _GEN_2555;
  reg  outputMemBlock_504;
  reg [31:0] _GEN_2556;
  reg  outputMemBlock_505;
  reg [31:0] _GEN_2557;
  reg  outputMemBlock_506;
  reg [31:0] _GEN_2558;
  reg  outputMemBlock_507;
  reg [31:0] _GEN_2559;
  reg  outputMemBlock_508;
  reg [31:0] _GEN_2560;
  reg  outputMemBlock_509;
  reg [31:0] _GEN_2561;
  reg  outputMemBlock_510;
  reg [31:0] _GEN_2562;
  reg  outputMemBlock_511;
  reg [31:0] _GEN_2563;
  reg [9:0] outputBits;
  reg [31:0] _GEN_2564;
  wire  nextBitValid;
  wire  nextBit;
  wire  inputAdvance;
  wire  _T_1579;
  wire  _T_1581;
  wire  _T_1582;
  wire [10:0] _T_1584;
  wire [9:0] _T_1585;
  wire [9:0] _GEN_513;
  wire  _GEN_514;
  wire  _GEN_515;
  wire  _GEN_516;
  wire  _GEN_517;
  wire  _GEN_518;
  wire  _GEN_519;
  wire  _GEN_520;
  wire  _GEN_521;
  wire  _GEN_522;
  wire  _GEN_523;
  wire  _GEN_524;
  wire  _GEN_525;
  wire  _GEN_526;
  wire  _GEN_527;
  wire  _GEN_528;
  wire  _GEN_529;
  wire  _GEN_530;
  wire  _GEN_531;
  wire  _GEN_532;
  wire  _GEN_533;
  wire  _GEN_534;
  wire  _GEN_535;
  wire  _GEN_536;
  wire  _GEN_537;
  wire  _GEN_538;
  wire  _GEN_539;
  wire  _GEN_540;
  wire  _GEN_541;
  wire  _GEN_542;
  wire  _GEN_543;
  wire  _GEN_544;
  wire  _GEN_545;
  wire  _GEN_546;
  wire  _GEN_547;
  wire  _GEN_548;
  wire  _GEN_549;
  wire  _GEN_550;
  wire  _GEN_551;
  wire  _GEN_552;
  wire  _GEN_553;
  wire  _GEN_554;
  wire  _GEN_555;
  wire  _GEN_556;
  wire  _GEN_557;
  wire  _GEN_558;
  wire  _GEN_559;
  wire  _GEN_560;
  wire  _GEN_561;
  wire  _GEN_562;
  wire  _GEN_563;
  wire  _GEN_564;
  wire  _GEN_565;
  wire  _GEN_566;
  wire  _GEN_567;
  wire  _GEN_568;
  wire  _GEN_569;
  wire  _GEN_570;
  wire  _GEN_571;
  wire  _GEN_572;
  wire  _GEN_573;
  wire  _GEN_574;
  wire  _GEN_575;
  wire  _GEN_576;
  wire  _GEN_577;
  wire  _GEN_578;
  wire  _GEN_579;
  wire  _GEN_580;
  wire  _GEN_581;
  wire  _GEN_582;
  wire  _GEN_583;
  wire  _GEN_584;
  wire  _GEN_585;
  wire  _GEN_586;
  wire  _GEN_587;
  wire  _GEN_588;
  wire  _GEN_589;
  wire  _GEN_590;
  wire  _GEN_591;
  wire  _GEN_592;
  wire  _GEN_593;
  wire  _GEN_594;
  wire  _GEN_595;
  wire  _GEN_596;
  wire  _GEN_597;
  wire  _GEN_598;
  wire  _GEN_599;
  wire  _GEN_600;
  wire  _GEN_601;
  wire  _GEN_602;
  wire  _GEN_603;
  wire  _GEN_604;
  wire  _GEN_605;
  wire  _GEN_606;
  wire  _GEN_607;
  wire  _GEN_608;
  wire  _GEN_609;
  wire  _GEN_610;
  wire  _GEN_611;
  wire  _GEN_612;
  wire  _GEN_613;
  wire  _GEN_614;
  wire  _GEN_615;
  wire  _GEN_616;
  wire  _GEN_617;
  wire  _GEN_618;
  wire  _GEN_619;
  wire  _GEN_620;
  wire  _GEN_621;
  wire  _GEN_622;
  wire  _GEN_623;
  wire  _GEN_624;
  wire  _GEN_625;
  wire  _GEN_626;
  wire  _GEN_627;
  wire  _GEN_628;
  wire  _GEN_629;
  wire  _GEN_630;
  wire  _GEN_631;
  wire  _GEN_632;
  wire  _GEN_633;
  wire  _GEN_634;
  wire  _GEN_635;
  wire  _GEN_636;
  wire  _GEN_637;
  wire  _GEN_638;
  wire  _GEN_639;
  wire  _GEN_640;
  wire  _GEN_641;
  wire  _GEN_642;
  wire  _GEN_643;
  wire  _GEN_644;
  wire  _GEN_645;
  wire  _GEN_646;
  wire  _GEN_647;
  wire  _GEN_648;
  wire  _GEN_649;
  wire  _GEN_650;
  wire  _GEN_651;
  wire  _GEN_652;
  wire  _GEN_653;
  wire  _GEN_654;
  wire  _GEN_655;
  wire  _GEN_656;
  wire  _GEN_657;
  wire  _GEN_658;
  wire  _GEN_659;
  wire  _GEN_660;
  wire  _GEN_661;
  wire  _GEN_662;
  wire  _GEN_663;
  wire  _GEN_664;
  wire  _GEN_665;
  wire  _GEN_666;
  wire  _GEN_667;
  wire  _GEN_668;
  wire  _GEN_669;
  wire  _GEN_670;
  wire  _GEN_671;
  wire  _GEN_672;
  wire  _GEN_673;
  wire  _GEN_674;
  wire  _GEN_675;
  wire  _GEN_676;
  wire  _GEN_677;
  wire  _GEN_678;
  wire  _GEN_679;
  wire  _GEN_680;
  wire  _GEN_681;
  wire  _GEN_682;
  wire  _GEN_683;
  wire  _GEN_684;
  wire  _GEN_685;
  wire  _GEN_686;
  wire  _GEN_687;
  wire  _GEN_688;
  wire  _GEN_689;
  wire  _GEN_690;
  wire  _GEN_691;
  wire  _GEN_692;
  wire  _GEN_693;
  wire  _GEN_694;
  wire  _GEN_695;
  wire  _GEN_696;
  wire  _GEN_697;
  wire  _GEN_698;
  wire  _GEN_699;
  wire  _GEN_700;
  wire  _GEN_701;
  wire  _GEN_702;
  wire  _GEN_703;
  wire  _GEN_704;
  wire  _GEN_705;
  wire  _GEN_706;
  wire  _GEN_707;
  wire  _GEN_708;
  wire  _GEN_709;
  wire  _GEN_710;
  wire  _GEN_711;
  wire  _GEN_712;
  wire  _GEN_713;
  wire  _GEN_714;
  wire  _GEN_715;
  wire  _GEN_716;
  wire  _GEN_717;
  wire  _GEN_718;
  wire  _GEN_719;
  wire  _GEN_720;
  wire  _GEN_721;
  wire  _GEN_722;
  wire  _GEN_723;
  wire  _GEN_724;
  wire  _GEN_725;
  wire  _GEN_726;
  wire  _GEN_727;
  wire  _GEN_728;
  wire  _GEN_729;
  wire  _GEN_730;
  wire  _GEN_731;
  wire  _GEN_732;
  wire  _GEN_733;
  wire  _GEN_734;
  wire  _GEN_735;
  wire  _GEN_736;
  wire  _GEN_737;
  wire  _GEN_738;
  wire  _GEN_739;
  wire  _GEN_740;
  wire  _GEN_741;
  wire  _GEN_742;
  wire  _GEN_743;
  wire  _GEN_744;
  wire  _GEN_745;
  wire  _GEN_746;
  wire  _GEN_747;
  wire  _GEN_748;
  wire  _GEN_749;
  wire  _GEN_750;
  wire  _GEN_751;
  wire  _GEN_752;
  wire  _GEN_753;
  wire  _GEN_754;
  wire  _GEN_755;
  wire  _GEN_756;
  wire  _GEN_757;
  wire  _GEN_758;
  wire  _GEN_759;
  wire  _GEN_760;
  wire  _GEN_761;
  wire  _GEN_762;
  wire  _GEN_763;
  wire  _GEN_764;
  wire  _GEN_765;
  wire  _GEN_766;
  wire  _GEN_767;
  wire  _GEN_768;
  wire  _GEN_769;
  wire  _GEN_770;
  wire  _GEN_771;
  wire  _GEN_772;
  wire  _GEN_773;
  wire  _GEN_774;
  wire  _GEN_775;
  wire  _GEN_776;
  wire  _GEN_777;
  wire  _GEN_778;
  wire  _GEN_779;
  wire  _GEN_780;
  wire  _GEN_781;
  wire  _GEN_782;
  wire  _GEN_783;
  wire  _GEN_784;
  wire  _GEN_785;
  wire  _GEN_786;
  wire  _GEN_787;
  wire  _GEN_788;
  wire  _GEN_789;
  wire  _GEN_790;
  wire  _GEN_791;
  wire  _GEN_792;
  wire  _GEN_793;
  wire  _GEN_794;
  wire  _GEN_795;
  wire  _GEN_796;
  wire  _GEN_797;
  wire  _GEN_798;
  wire  _GEN_799;
  wire  _GEN_800;
  wire  _GEN_801;
  wire  _GEN_802;
  wire  _GEN_803;
  wire  _GEN_804;
  wire  _GEN_805;
  wire  _GEN_806;
  wire  _GEN_807;
  wire  _GEN_808;
  wire  _GEN_809;
  wire  _GEN_810;
  wire  _GEN_811;
  wire  _GEN_812;
  wire  _GEN_813;
  wire  _GEN_814;
  wire  _GEN_815;
  wire  _GEN_816;
  wire  _GEN_817;
  wire  _GEN_818;
  wire  _GEN_819;
  wire  _GEN_820;
  wire  _GEN_821;
  wire  _GEN_822;
  wire  _GEN_823;
  wire  _GEN_824;
  wire  _GEN_825;
  wire  _GEN_826;
  wire  _GEN_827;
  wire  _GEN_828;
  wire  _GEN_829;
  wire  _GEN_830;
  wire  _GEN_831;
  wire  _GEN_832;
  wire  _GEN_833;
  wire  _GEN_834;
  wire  _GEN_835;
  wire  _GEN_836;
  wire  _GEN_837;
  wire  _GEN_838;
  wire  _GEN_839;
  wire  _GEN_840;
  wire  _GEN_841;
  wire  _GEN_842;
  wire  _GEN_843;
  wire  _GEN_844;
  wire  _GEN_845;
  wire  _GEN_846;
  wire  _GEN_847;
  wire  _GEN_848;
  wire  _GEN_849;
  wire  _GEN_850;
  wire  _GEN_851;
  wire  _GEN_852;
  wire  _GEN_853;
  wire  _GEN_854;
  wire  _GEN_855;
  wire  _GEN_856;
  wire  _GEN_857;
  wire  _GEN_858;
  wire  _GEN_859;
  wire  _GEN_860;
  wire  _GEN_861;
  wire  _GEN_862;
  wire  _GEN_863;
  wire  _GEN_864;
  wire  _GEN_865;
  wire  _GEN_866;
  wire  _GEN_867;
  wire  _GEN_868;
  wire  _GEN_869;
  wire  _GEN_870;
  wire  _GEN_871;
  wire  _GEN_872;
  wire  _GEN_873;
  wire  _GEN_874;
  wire  _GEN_875;
  wire  _GEN_876;
  wire  _GEN_877;
  wire  _GEN_878;
  wire  _GEN_879;
  wire  _GEN_880;
  wire  _GEN_881;
  wire  _GEN_882;
  wire  _GEN_883;
  wire  _GEN_884;
  wire  _GEN_885;
  wire  _GEN_886;
  wire  _GEN_887;
  wire  _GEN_888;
  wire  _GEN_889;
  wire  _GEN_890;
  wire  _GEN_891;
  wire  _GEN_892;
  wire  _GEN_893;
  wire  _GEN_894;
  wire  _GEN_895;
  wire  _GEN_896;
  wire  _GEN_897;
  wire  _GEN_898;
  wire  _GEN_899;
  wire  _GEN_900;
  wire  _GEN_901;
  wire  _GEN_902;
  wire  _GEN_903;
  wire  _GEN_904;
  wire  _GEN_905;
  wire  _GEN_906;
  wire  _GEN_907;
  wire  _GEN_908;
  wire  _GEN_909;
  wire  _GEN_910;
  wire  _GEN_911;
  wire  _GEN_912;
  wire  _GEN_913;
  wire  _GEN_914;
  wire  _GEN_915;
  wire  _GEN_916;
  wire  _GEN_917;
  wire  _GEN_918;
  wire  _GEN_919;
  wire  _GEN_920;
  wire  _GEN_921;
  wire  _GEN_922;
  wire  _GEN_923;
  wire  _GEN_924;
  wire  _GEN_925;
  wire  _GEN_926;
  wire  _GEN_927;
  wire  _GEN_928;
  wire  _GEN_929;
  wire  _GEN_930;
  wire  _GEN_931;
  wire  _GEN_932;
  wire  _GEN_933;
  wire  _GEN_934;
  wire  _GEN_935;
  wire  _GEN_936;
  wire  _GEN_937;
  wire  _GEN_938;
  wire  _GEN_939;
  wire  _GEN_940;
  wire  _GEN_941;
  wire  _GEN_942;
  wire  _GEN_943;
  wire  _GEN_944;
  wire  _GEN_945;
  wire  _GEN_946;
  wire  _GEN_947;
  wire  _GEN_948;
  wire  _GEN_949;
  wire  _GEN_950;
  wire  _GEN_951;
  wire  _GEN_952;
  wire  _GEN_953;
  wire  _GEN_954;
  wire  _GEN_955;
  wire  _GEN_956;
  wire  _GEN_957;
  wire  _GEN_958;
  wire  _GEN_959;
  wire  _GEN_960;
  wire  _GEN_961;
  wire  _GEN_962;
  wire  _GEN_963;
  wire  _GEN_964;
  wire  _GEN_965;
  wire  _GEN_966;
  wire  _GEN_967;
  wire  _GEN_968;
  wire  _GEN_969;
  wire  _GEN_970;
  wire  _GEN_971;
  wire  _GEN_972;
  wire  _GEN_973;
  wire  _GEN_974;
  wire  _GEN_975;
  wire  _GEN_976;
  wire  _GEN_977;
  wire  _GEN_978;
  wire  _GEN_979;
  wire  _GEN_980;
  wire  _GEN_981;
  wire  _GEN_982;
  wire  _GEN_983;
  wire  _GEN_984;
  wire  _GEN_985;
  wire  _GEN_986;
  wire  _GEN_987;
  wire  _GEN_988;
  wire  _GEN_989;
  wire  _GEN_990;
  wire  _GEN_991;
  wire  _GEN_992;
  wire  _GEN_993;
  wire  _GEN_994;
  wire  _GEN_995;
  wire  _GEN_996;
  wire  _GEN_997;
  wire  _GEN_998;
  wire  _GEN_999;
  wire  _GEN_1000;
  wire  _GEN_1001;
  wire  _GEN_1002;
  wire  _GEN_1003;
  wire  _GEN_1004;
  wire  _GEN_1005;
  wire  _GEN_1006;
  wire  _GEN_1007;
  wire  _GEN_1008;
  wire  _GEN_1009;
  wire  _GEN_1010;
  wire  _GEN_1011;
  wire  _GEN_1012;
  wire  _GEN_1013;
  wire  _GEN_1014;
  wire  _GEN_1015;
  wire  _GEN_1016;
  wire  _GEN_1017;
  wire  _GEN_1018;
  wire  _GEN_1019;
  wire  _GEN_1020;
  wire  _GEN_1021;
  wire  _GEN_1022;
  wire  _GEN_1023;
  wire  _GEN_1024;
  wire [10:0] _T_1587;
  wire [9:0] _T_1588;
  wire  _GEN_1025;
  wire  _GEN_1026;
  wire  _GEN_1027;
  wire  _GEN_1028;
  wire  _GEN_1029;
  wire  _GEN_1030;
  wire  _GEN_1031;
  wire  _GEN_1032;
  wire  _GEN_1033;
  wire  _GEN_1034;
  wire  _GEN_1035;
  wire  _GEN_1036;
  wire  _GEN_1037;
  wire  _GEN_1038;
  wire  _GEN_1039;
  wire  _GEN_1040;
  wire  _GEN_1041;
  wire  _GEN_1042;
  wire  _GEN_1043;
  wire  _GEN_1044;
  wire  _GEN_1045;
  wire  _GEN_1046;
  wire  _GEN_1047;
  wire  _GEN_1048;
  wire  _GEN_1049;
  wire  _GEN_1050;
  wire  _GEN_1051;
  wire  _GEN_1052;
  wire  _GEN_1053;
  wire  _GEN_1054;
  wire  _GEN_1055;
  wire  _GEN_1056;
  wire  _GEN_1057;
  wire  _GEN_1058;
  wire  _GEN_1059;
  wire  _GEN_1060;
  wire  _GEN_1061;
  wire  _GEN_1062;
  wire  _GEN_1063;
  wire  _GEN_1064;
  wire  _GEN_1065;
  wire  _GEN_1066;
  wire  _GEN_1067;
  wire  _GEN_1068;
  wire  _GEN_1069;
  wire  _GEN_1070;
  wire  _GEN_1071;
  wire  _GEN_1072;
  wire  _GEN_1073;
  wire  _GEN_1074;
  wire  _GEN_1075;
  wire  _GEN_1076;
  wire  _GEN_1077;
  wire  _GEN_1078;
  wire  _GEN_1079;
  wire  _GEN_1080;
  wire  _GEN_1081;
  wire  _GEN_1082;
  wire  _GEN_1083;
  wire  _GEN_1084;
  wire  _GEN_1085;
  wire  _GEN_1086;
  wire  _GEN_1087;
  wire  _GEN_1088;
  wire  _GEN_1089;
  wire  _GEN_1090;
  wire  _GEN_1091;
  wire  _GEN_1092;
  wire  _GEN_1093;
  wire  _GEN_1094;
  wire  _GEN_1095;
  wire  _GEN_1096;
  wire  _GEN_1097;
  wire  _GEN_1098;
  wire  _GEN_1099;
  wire  _GEN_1100;
  wire  _GEN_1101;
  wire  _GEN_1102;
  wire  _GEN_1103;
  wire  _GEN_1104;
  wire  _GEN_1105;
  wire  _GEN_1106;
  wire  _GEN_1107;
  wire  _GEN_1108;
  wire  _GEN_1109;
  wire  _GEN_1110;
  wire  _GEN_1111;
  wire  _GEN_1112;
  wire  _GEN_1113;
  wire  _GEN_1114;
  wire  _GEN_1115;
  wire  _GEN_1116;
  wire  _GEN_1117;
  wire  _GEN_1118;
  wire  _GEN_1119;
  wire  _GEN_1120;
  wire  _GEN_1121;
  wire  _GEN_1122;
  wire  _GEN_1123;
  wire  _GEN_1124;
  wire  _GEN_1125;
  wire  _GEN_1126;
  wire  _GEN_1127;
  wire  _GEN_1128;
  wire  _GEN_1129;
  wire  _GEN_1130;
  wire  _GEN_1131;
  wire  _GEN_1132;
  wire  _GEN_1133;
  wire  _GEN_1134;
  wire  _GEN_1135;
  wire  _GEN_1136;
  wire  _GEN_1137;
  wire  _GEN_1138;
  wire  _GEN_1139;
  wire  _GEN_1140;
  wire  _GEN_1141;
  wire  _GEN_1142;
  wire  _GEN_1143;
  wire  _GEN_1144;
  wire  _GEN_1145;
  wire  _GEN_1146;
  wire  _GEN_1147;
  wire  _GEN_1148;
  wire  _GEN_1149;
  wire  _GEN_1150;
  wire  _GEN_1151;
  wire  _GEN_1152;
  wire  _GEN_1153;
  wire  _GEN_1154;
  wire  _GEN_1155;
  wire  _GEN_1156;
  wire  _GEN_1157;
  wire  _GEN_1158;
  wire  _GEN_1159;
  wire  _GEN_1160;
  wire  _GEN_1161;
  wire  _GEN_1162;
  wire  _GEN_1163;
  wire  _GEN_1164;
  wire  _GEN_1165;
  wire  _GEN_1166;
  wire  _GEN_1167;
  wire  _GEN_1168;
  wire  _GEN_1169;
  wire  _GEN_1170;
  wire  _GEN_1171;
  wire  _GEN_1172;
  wire  _GEN_1173;
  wire  _GEN_1174;
  wire  _GEN_1175;
  wire  _GEN_1176;
  wire  _GEN_1177;
  wire  _GEN_1178;
  wire  _GEN_1179;
  wire  _GEN_1180;
  wire  _GEN_1181;
  wire  _GEN_1182;
  wire  _GEN_1183;
  wire  _GEN_1184;
  wire  _GEN_1185;
  wire  _GEN_1186;
  wire  _GEN_1187;
  wire  _GEN_1188;
  wire  _GEN_1189;
  wire  _GEN_1190;
  wire  _GEN_1191;
  wire  _GEN_1192;
  wire  _GEN_1193;
  wire  _GEN_1194;
  wire  _GEN_1195;
  wire  _GEN_1196;
  wire  _GEN_1197;
  wire  _GEN_1198;
  wire  _GEN_1199;
  wire  _GEN_1200;
  wire  _GEN_1201;
  wire  _GEN_1202;
  wire  _GEN_1203;
  wire  _GEN_1204;
  wire  _GEN_1205;
  wire  _GEN_1206;
  wire  _GEN_1207;
  wire  _GEN_1208;
  wire  _GEN_1209;
  wire  _GEN_1210;
  wire  _GEN_1211;
  wire  _GEN_1212;
  wire  _GEN_1213;
  wire  _GEN_1214;
  wire  _GEN_1215;
  wire  _GEN_1216;
  wire  _GEN_1217;
  wire  _GEN_1218;
  wire  _GEN_1219;
  wire  _GEN_1220;
  wire  _GEN_1221;
  wire  _GEN_1222;
  wire  _GEN_1223;
  wire  _GEN_1224;
  wire  _GEN_1225;
  wire  _GEN_1226;
  wire  _GEN_1227;
  wire  _GEN_1228;
  wire  _GEN_1229;
  wire  _GEN_1230;
  wire  _GEN_1231;
  wire  _GEN_1232;
  wire  _GEN_1233;
  wire  _GEN_1234;
  wire  _GEN_1235;
  wire  _GEN_1236;
  wire  _GEN_1237;
  wire  _GEN_1238;
  wire  _GEN_1239;
  wire  _GEN_1240;
  wire  _GEN_1241;
  wire  _GEN_1242;
  wire  _GEN_1243;
  wire  _GEN_1244;
  wire  _GEN_1245;
  wire  _GEN_1246;
  wire  _GEN_1247;
  wire  _GEN_1248;
  wire  _GEN_1249;
  wire  _GEN_1250;
  wire  _GEN_1251;
  wire  _GEN_1252;
  wire  _GEN_1253;
  wire  _GEN_1254;
  wire  _GEN_1255;
  wire  _GEN_1256;
  wire  _GEN_1257;
  wire  _GEN_1258;
  wire  _GEN_1259;
  wire  _GEN_1260;
  wire  _GEN_1261;
  wire  _GEN_1262;
  wire  _GEN_1263;
  wire  _GEN_1264;
  wire  _GEN_1265;
  wire  _GEN_1266;
  wire  _GEN_1267;
  wire  _GEN_1268;
  wire  _GEN_1269;
  wire  _GEN_1270;
  wire  _GEN_1271;
  wire  _GEN_1272;
  wire  _GEN_1273;
  wire  _GEN_1274;
  wire  _GEN_1275;
  wire  _GEN_1276;
  wire  _GEN_1277;
  wire  _GEN_1278;
  wire  _GEN_1279;
  wire  _GEN_1280;
  wire  _GEN_1281;
  wire  _GEN_1282;
  wire  _GEN_1283;
  wire  _GEN_1284;
  wire  _GEN_1285;
  wire  _GEN_1286;
  wire  _GEN_1287;
  wire  _GEN_1288;
  wire  _GEN_1289;
  wire  _GEN_1290;
  wire  _GEN_1291;
  wire  _GEN_1292;
  wire  _GEN_1293;
  wire  _GEN_1294;
  wire  _GEN_1295;
  wire  _GEN_1296;
  wire  _GEN_1297;
  wire  _GEN_1298;
  wire  _GEN_1299;
  wire  _GEN_1300;
  wire  _GEN_1301;
  wire  _GEN_1302;
  wire  _GEN_1303;
  wire  _GEN_1304;
  wire  _GEN_1305;
  wire  _GEN_1306;
  wire  _GEN_1307;
  wire  _GEN_1308;
  wire  _GEN_1309;
  wire  _GEN_1310;
  wire  _GEN_1311;
  wire  _GEN_1312;
  wire  _GEN_1313;
  wire  _GEN_1314;
  wire  _GEN_1315;
  wire  _GEN_1316;
  wire  _GEN_1317;
  wire  _GEN_1318;
  wire  _GEN_1319;
  wire  _GEN_1320;
  wire  _GEN_1321;
  wire  _GEN_1322;
  wire  _GEN_1323;
  wire  _GEN_1324;
  wire  _GEN_1325;
  wire  _GEN_1326;
  wire  _GEN_1327;
  wire  _GEN_1328;
  wire  _GEN_1329;
  wire  _GEN_1330;
  wire  _GEN_1331;
  wire  _GEN_1332;
  wire  _GEN_1333;
  wire  _GEN_1334;
  wire  _GEN_1335;
  wire  _GEN_1336;
  wire  _GEN_1337;
  wire  _GEN_1338;
  wire  _GEN_1339;
  wire  _GEN_1340;
  wire  _GEN_1341;
  wire  _GEN_1342;
  wire  _GEN_1343;
  wire  _GEN_1344;
  wire  _GEN_1345;
  wire  _GEN_1346;
  wire  _GEN_1347;
  wire  _GEN_1348;
  wire  _GEN_1349;
  wire  _GEN_1350;
  wire  _GEN_1351;
  wire  _GEN_1352;
  wire  _GEN_1353;
  wire  _GEN_1354;
  wire  _GEN_1355;
  wire  _GEN_1356;
  wire  _GEN_1357;
  wire  _GEN_1358;
  wire  _GEN_1359;
  wire  _GEN_1360;
  wire  _GEN_1361;
  wire  _GEN_1362;
  wire  _GEN_1363;
  wire  _GEN_1364;
  wire  _GEN_1365;
  wire  _GEN_1366;
  wire  _GEN_1367;
  wire  _GEN_1368;
  wire  _GEN_1369;
  wire  _GEN_1370;
  wire  _GEN_1371;
  wire  _GEN_1372;
  wire  _GEN_1373;
  wire  _GEN_1374;
  wire  _GEN_1375;
  wire  _GEN_1376;
  wire  _GEN_1377;
  wire  _GEN_1378;
  wire  _GEN_1379;
  wire  _GEN_1380;
  wire  _GEN_1381;
  wire  _GEN_1382;
  wire  _GEN_1383;
  wire  _GEN_1384;
  wire  _GEN_1385;
  wire  _GEN_1386;
  wire  _GEN_1387;
  wire  _GEN_1388;
  wire  _GEN_1389;
  wire  _GEN_1390;
  wire  _GEN_1391;
  wire  _GEN_1392;
  wire  _GEN_1393;
  wire  _GEN_1394;
  wire  _GEN_1395;
  wire  _GEN_1396;
  wire  _GEN_1397;
  wire  _GEN_1398;
  wire  _GEN_1399;
  wire  _GEN_1400;
  wire  _GEN_1401;
  wire  _GEN_1402;
  wire  _GEN_1403;
  wire  _GEN_1404;
  wire  _GEN_1405;
  wire  _GEN_1406;
  wire  _GEN_1407;
  wire  _GEN_1408;
  wire  _GEN_1409;
  wire  _GEN_1410;
  wire  _GEN_1411;
  wire  _GEN_1412;
  wire  _GEN_1413;
  wire  _GEN_1414;
  wire  _GEN_1415;
  wire  _GEN_1416;
  wire  _GEN_1417;
  wire  _GEN_1418;
  wire  _GEN_1419;
  wire  _GEN_1420;
  wire  _GEN_1421;
  wire  _GEN_1422;
  wire  _GEN_1423;
  wire  _GEN_1424;
  wire  _GEN_1425;
  wire  _GEN_1426;
  wire  _GEN_1427;
  wire  _GEN_1428;
  wire  _GEN_1429;
  wire  _GEN_1430;
  wire  _GEN_1431;
  wire  _GEN_1432;
  wire  _GEN_1433;
  wire  _GEN_1434;
  wire  _GEN_1435;
  wire  _GEN_1436;
  wire  _GEN_1437;
  wire  _GEN_1438;
  wire  _GEN_1439;
  wire  _GEN_1440;
  wire  _GEN_1441;
  wire  _GEN_1442;
  wire  _GEN_1443;
  wire  _GEN_1444;
  wire  _GEN_1445;
  wire  _GEN_1446;
  wire  _GEN_1447;
  wire  _GEN_1448;
  wire  _GEN_1449;
  wire  _GEN_1450;
  wire  _GEN_1451;
  wire  _GEN_1452;
  wire  _GEN_1453;
  wire  _GEN_1454;
  wire  _GEN_1455;
  wire  _GEN_1456;
  wire  _GEN_1457;
  wire  _GEN_1458;
  wire  _GEN_1459;
  wire  _GEN_1460;
  wire  _GEN_1461;
  wire  _GEN_1462;
  wire  _GEN_1463;
  wire  _GEN_1464;
  wire  _GEN_1465;
  wire  _GEN_1466;
  wire  _GEN_1467;
  wire  _GEN_1468;
  wire  _GEN_1469;
  wire  _GEN_1470;
  wire  _GEN_1471;
  wire  _GEN_1472;
  wire  _GEN_1473;
  wire  _GEN_1474;
  wire  _GEN_1475;
  wire  _GEN_1476;
  wire  _GEN_1477;
  wire  _GEN_1478;
  wire  _GEN_1479;
  wire  _GEN_1480;
  wire  _GEN_1481;
  wire  _GEN_1482;
  wire  _GEN_1483;
  wire  _GEN_1484;
  wire  _GEN_1485;
  wire  _GEN_1486;
  wire  _GEN_1487;
  wire  _GEN_1488;
  wire  _GEN_1489;
  wire  _GEN_1490;
  wire  _GEN_1491;
  wire  _GEN_1492;
  wire  _GEN_1493;
  wire  _GEN_1494;
  wire  _GEN_1495;
  wire  _GEN_1496;
  wire  _GEN_1497;
  wire  _GEN_1498;
  wire  _GEN_1499;
  wire  _GEN_1500;
  wire  _GEN_1501;
  wire  _GEN_1502;
  wire  _GEN_1503;
  wire  _GEN_1504;
  wire  _GEN_1505;
  wire  _GEN_1506;
  wire  _GEN_1507;
  wire  _GEN_1508;
  wire  _GEN_1509;
  wire  _GEN_1510;
  wire  _GEN_1511;
  wire  _GEN_1512;
  wire  _GEN_1513;
  wire  _GEN_1514;
  wire  _GEN_1515;
  wire  _GEN_1516;
  wire  _GEN_1517;
  wire  _GEN_1518;
  wire  _GEN_1519;
  wire  _GEN_1520;
  wire  _GEN_1521;
  wire  _GEN_1522;
  wire  _GEN_1523;
  wire  _GEN_1524;
  wire  _GEN_1525;
  wire  _GEN_1526;
  wire  _GEN_1527;
  wire  _GEN_1528;
  wire  _GEN_1529;
  wire  _GEN_1530;
  wire  _GEN_1531;
  wire  _GEN_1532;
  wire  _GEN_1533;
  wire  _GEN_1534;
  wire  _GEN_1535;
  wire  _GEN_1536;
  wire [9:0] _GEN_1537;
  wire  _T_1590;
  wire  _T_1593;
  wire  _T_1595;
  wire  _T_1596;
  wire  _T_1597;
  wire [1:0] _T_1598;
  wire [1:0] _T_1599;
  wire [3:0] _T_1600;
  wire [1:0] _T_1601;
  wire [1:0] _T_1602;
  wire [3:0] _T_1603;
  wire [7:0] _T_1604;
  wire [1:0] _T_1605;
  wire [1:0] _T_1606;
  wire [3:0] _T_1607;
  wire [1:0] _T_1608;
  wire [1:0] _T_1609;
  wire [3:0] _T_1610;
  wire [7:0] _T_1611;
  wire [15:0] _T_1612;
  wire [1:0] _T_1613;
  wire [1:0] _T_1614;
  wire [3:0] _T_1615;
  wire [1:0] _T_1616;
  wire [1:0] _T_1617;
  wire [3:0] _T_1618;
  wire [7:0] _T_1619;
  wire [1:0] _T_1620;
  wire [1:0] _T_1621;
  wire [3:0] _T_1622;
  wire [1:0] _T_1623;
  wire [1:0] _T_1624;
  wire [3:0] _T_1625;
  wire [7:0] _T_1626;
  wire [15:0] _T_1627;
  wire [31:0] _T_1628;
  wire [1:0] _T_1629;
  wire [1:0] _T_1630;
  wire [3:0] _T_1631;
  wire [1:0] _T_1632;
  wire [1:0] _T_1633;
  wire [3:0] _T_1634;
  wire [7:0] _T_1635;
  wire [1:0] _T_1636;
  wire [1:0] _T_1637;
  wire [3:0] _T_1638;
  wire [1:0] _T_1639;
  wire [1:0] _T_1640;
  wire [3:0] _T_1641;
  wire [7:0] _T_1642;
  wire [15:0] _T_1643;
  wire [1:0] _T_1644;
  wire [1:0] _T_1645;
  wire [3:0] _T_1646;
  wire [1:0] _T_1647;
  wire [1:0] _T_1648;
  wire [3:0] _T_1649;
  wire [7:0] _T_1650;
  wire [1:0] _T_1651;
  wire [1:0] _T_1652;
  wire [3:0] _T_1653;
  wire [1:0] _T_1654;
  wire [1:0] _T_1655;
  wire [3:0] _T_1656;
  wire [7:0] _T_1657;
  wire [15:0] _T_1658;
  wire [31:0] _T_1659;
  wire [63:0] _T_1660;
  wire [1:0] _T_1661;
  wire [1:0] _T_1662;
  wire [3:0] _T_1663;
  wire [1:0] _T_1664;
  wire [1:0] _T_1665;
  wire [3:0] _T_1666;
  wire [7:0] _T_1667;
  wire [1:0] _T_1668;
  wire [1:0] _T_1669;
  wire [3:0] _T_1670;
  wire [1:0] _T_1671;
  wire [1:0] _T_1672;
  wire [3:0] _T_1673;
  wire [7:0] _T_1674;
  wire [15:0] _T_1675;
  wire [1:0] _T_1676;
  wire [1:0] _T_1677;
  wire [3:0] _T_1678;
  wire [1:0] _T_1679;
  wire [1:0] _T_1680;
  wire [3:0] _T_1681;
  wire [7:0] _T_1682;
  wire [1:0] _T_1683;
  wire [1:0] _T_1684;
  wire [3:0] _T_1685;
  wire [1:0] _T_1686;
  wire [1:0] _T_1687;
  wire [3:0] _T_1688;
  wire [7:0] _T_1689;
  wire [15:0] _T_1690;
  wire [31:0] _T_1691;
  wire [1:0] _T_1692;
  wire [1:0] _T_1693;
  wire [3:0] _T_1694;
  wire [1:0] _T_1695;
  wire [1:0] _T_1696;
  wire [3:0] _T_1697;
  wire [7:0] _T_1698;
  wire [1:0] _T_1699;
  wire [1:0] _T_1700;
  wire [3:0] _T_1701;
  wire [1:0] _T_1702;
  wire [1:0] _T_1703;
  wire [3:0] _T_1704;
  wire [7:0] _T_1705;
  wire [15:0] _T_1706;
  wire [1:0] _T_1707;
  wire [1:0] _T_1708;
  wire [3:0] _T_1709;
  wire [1:0] _T_1710;
  wire [1:0] _T_1711;
  wire [3:0] _T_1712;
  wire [7:0] _T_1713;
  wire [1:0] _T_1714;
  wire [1:0] _T_1715;
  wire [3:0] _T_1716;
  wire [1:0] _T_1717;
  wire [1:0] _T_1718;
  wire [3:0] _T_1719;
  wire [7:0] _T_1720;
  wire [15:0] _T_1721;
  wire [31:0] _T_1722;
  wire [63:0] _T_1723;
  wire [127:0] _T_1724;
  wire [1:0] _T_1725;
  wire [1:0] _T_1726;
  wire [3:0] _T_1727;
  wire [1:0] _T_1728;
  wire [1:0] _T_1729;
  wire [3:0] _T_1730;
  wire [7:0] _T_1731;
  wire [1:0] _T_1732;
  wire [1:0] _T_1733;
  wire [3:0] _T_1734;
  wire [1:0] _T_1735;
  wire [1:0] _T_1736;
  wire [3:0] _T_1737;
  wire [7:0] _T_1738;
  wire [15:0] _T_1739;
  wire [1:0] _T_1740;
  wire [1:0] _T_1741;
  wire [3:0] _T_1742;
  wire [1:0] _T_1743;
  wire [1:0] _T_1744;
  wire [3:0] _T_1745;
  wire [7:0] _T_1746;
  wire [1:0] _T_1747;
  wire [1:0] _T_1748;
  wire [3:0] _T_1749;
  wire [1:0] _T_1750;
  wire [1:0] _T_1751;
  wire [3:0] _T_1752;
  wire [7:0] _T_1753;
  wire [15:0] _T_1754;
  wire [31:0] _T_1755;
  wire [1:0] _T_1756;
  wire [1:0] _T_1757;
  wire [3:0] _T_1758;
  wire [1:0] _T_1759;
  wire [1:0] _T_1760;
  wire [3:0] _T_1761;
  wire [7:0] _T_1762;
  wire [1:0] _T_1763;
  wire [1:0] _T_1764;
  wire [3:0] _T_1765;
  wire [1:0] _T_1766;
  wire [1:0] _T_1767;
  wire [3:0] _T_1768;
  wire [7:0] _T_1769;
  wire [15:0] _T_1770;
  wire [1:0] _T_1771;
  wire [1:0] _T_1772;
  wire [3:0] _T_1773;
  wire [1:0] _T_1774;
  wire [1:0] _T_1775;
  wire [3:0] _T_1776;
  wire [7:0] _T_1777;
  wire [1:0] _T_1778;
  wire [1:0] _T_1779;
  wire [3:0] _T_1780;
  wire [1:0] _T_1781;
  wire [1:0] _T_1782;
  wire [3:0] _T_1783;
  wire [7:0] _T_1784;
  wire [15:0] _T_1785;
  wire [31:0] _T_1786;
  wire [63:0] _T_1787;
  wire [1:0] _T_1788;
  wire [1:0] _T_1789;
  wire [3:0] _T_1790;
  wire [1:0] _T_1791;
  wire [1:0] _T_1792;
  wire [3:0] _T_1793;
  wire [7:0] _T_1794;
  wire [1:0] _T_1795;
  wire [1:0] _T_1796;
  wire [3:0] _T_1797;
  wire [1:0] _T_1798;
  wire [1:0] _T_1799;
  wire [3:0] _T_1800;
  wire [7:0] _T_1801;
  wire [15:0] _T_1802;
  wire [1:0] _T_1803;
  wire [1:0] _T_1804;
  wire [3:0] _T_1805;
  wire [1:0] _T_1806;
  wire [1:0] _T_1807;
  wire [3:0] _T_1808;
  wire [7:0] _T_1809;
  wire [1:0] _T_1810;
  wire [1:0] _T_1811;
  wire [3:0] _T_1812;
  wire [1:0] _T_1813;
  wire [1:0] _T_1814;
  wire [3:0] _T_1815;
  wire [7:0] _T_1816;
  wire [15:0] _T_1817;
  wire [31:0] _T_1818;
  wire [1:0] _T_1819;
  wire [1:0] _T_1820;
  wire [3:0] _T_1821;
  wire [1:0] _T_1822;
  wire [1:0] _T_1823;
  wire [3:0] _T_1824;
  wire [7:0] _T_1825;
  wire [1:0] _T_1826;
  wire [1:0] _T_1827;
  wire [3:0] _T_1828;
  wire [1:0] _T_1829;
  wire [1:0] _T_1830;
  wire [3:0] _T_1831;
  wire [7:0] _T_1832;
  wire [15:0] _T_1833;
  wire [1:0] _T_1834;
  wire [1:0] _T_1835;
  wire [3:0] _T_1836;
  wire [1:0] _T_1837;
  wire [1:0] _T_1838;
  wire [3:0] _T_1839;
  wire [7:0] _T_1840;
  wire [1:0] _T_1841;
  wire [1:0] _T_1842;
  wire [3:0] _T_1843;
  wire [1:0] _T_1844;
  wire [1:0] _T_1845;
  wire [3:0] _T_1846;
  wire [7:0] _T_1847;
  wire [15:0] _T_1848;
  wire [31:0] _T_1849;
  wire [63:0] _T_1850;
  wire [127:0] _T_1851;
  wire [255:0] _T_1852;
  wire [1:0] _T_1853;
  wire [1:0] _T_1854;
  wire [3:0] _T_1855;
  wire [1:0] _T_1856;
  wire [1:0] _T_1857;
  wire [3:0] _T_1858;
  wire [7:0] _T_1859;
  wire [1:0] _T_1860;
  wire [1:0] _T_1861;
  wire [3:0] _T_1862;
  wire [1:0] _T_1863;
  wire [1:0] _T_1864;
  wire [3:0] _T_1865;
  wire [7:0] _T_1866;
  wire [15:0] _T_1867;
  wire [1:0] _T_1868;
  wire [1:0] _T_1869;
  wire [3:0] _T_1870;
  wire [1:0] _T_1871;
  wire [1:0] _T_1872;
  wire [3:0] _T_1873;
  wire [7:0] _T_1874;
  wire [1:0] _T_1875;
  wire [1:0] _T_1876;
  wire [3:0] _T_1877;
  wire [1:0] _T_1878;
  wire [1:0] _T_1879;
  wire [3:0] _T_1880;
  wire [7:0] _T_1881;
  wire [15:0] _T_1882;
  wire [31:0] _T_1883;
  wire [1:0] _T_1884;
  wire [1:0] _T_1885;
  wire [3:0] _T_1886;
  wire [1:0] _T_1887;
  wire [1:0] _T_1888;
  wire [3:0] _T_1889;
  wire [7:0] _T_1890;
  wire [1:0] _T_1891;
  wire [1:0] _T_1892;
  wire [3:0] _T_1893;
  wire [1:0] _T_1894;
  wire [1:0] _T_1895;
  wire [3:0] _T_1896;
  wire [7:0] _T_1897;
  wire [15:0] _T_1898;
  wire [1:0] _T_1899;
  wire [1:0] _T_1900;
  wire [3:0] _T_1901;
  wire [1:0] _T_1902;
  wire [1:0] _T_1903;
  wire [3:0] _T_1904;
  wire [7:0] _T_1905;
  wire [1:0] _T_1906;
  wire [1:0] _T_1907;
  wire [3:0] _T_1908;
  wire [1:0] _T_1909;
  wire [1:0] _T_1910;
  wire [3:0] _T_1911;
  wire [7:0] _T_1912;
  wire [15:0] _T_1913;
  wire [31:0] _T_1914;
  wire [63:0] _T_1915;
  wire [1:0] _T_1916;
  wire [1:0] _T_1917;
  wire [3:0] _T_1918;
  wire [1:0] _T_1919;
  wire [1:0] _T_1920;
  wire [3:0] _T_1921;
  wire [7:0] _T_1922;
  wire [1:0] _T_1923;
  wire [1:0] _T_1924;
  wire [3:0] _T_1925;
  wire [1:0] _T_1926;
  wire [1:0] _T_1927;
  wire [3:0] _T_1928;
  wire [7:0] _T_1929;
  wire [15:0] _T_1930;
  wire [1:0] _T_1931;
  wire [1:0] _T_1932;
  wire [3:0] _T_1933;
  wire [1:0] _T_1934;
  wire [1:0] _T_1935;
  wire [3:0] _T_1936;
  wire [7:0] _T_1937;
  wire [1:0] _T_1938;
  wire [1:0] _T_1939;
  wire [3:0] _T_1940;
  wire [1:0] _T_1941;
  wire [1:0] _T_1942;
  wire [3:0] _T_1943;
  wire [7:0] _T_1944;
  wire [15:0] _T_1945;
  wire [31:0] _T_1946;
  wire [1:0] _T_1947;
  wire [1:0] _T_1948;
  wire [3:0] _T_1949;
  wire [1:0] _T_1950;
  wire [1:0] _T_1951;
  wire [3:0] _T_1952;
  wire [7:0] _T_1953;
  wire [1:0] _T_1954;
  wire [1:0] _T_1955;
  wire [3:0] _T_1956;
  wire [1:0] _T_1957;
  wire [1:0] _T_1958;
  wire [3:0] _T_1959;
  wire [7:0] _T_1960;
  wire [15:0] _T_1961;
  wire [1:0] _T_1962;
  wire [1:0] _T_1963;
  wire [3:0] _T_1964;
  wire [1:0] _T_1965;
  wire [1:0] _T_1966;
  wire [3:0] _T_1967;
  wire [7:0] _T_1968;
  wire [1:0] _T_1969;
  wire [1:0] _T_1970;
  wire [3:0] _T_1971;
  wire [1:0] _T_1972;
  wire [1:0] _T_1973;
  wire [3:0] _T_1974;
  wire [7:0] _T_1975;
  wire [15:0] _T_1976;
  wire [31:0] _T_1977;
  wire [63:0] _T_1978;
  wire [127:0] _T_1979;
  wire [1:0] _T_1980;
  wire [1:0] _T_1981;
  wire [3:0] _T_1982;
  wire [1:0] _T_1983;
  wire [1:0] _T_1984;
  wire [3:0] _T_1985;
  wire [7:0] _T_1986;
  wire [1:0] _T_1987;
  wire [1:0] _T_1988;
  wire [3:0] _T_1989;
  wire [1:0] _T_1990;
  wire [1:0] _T_1991;
  wire [3:0] _T_1992;
  wire [7:0] _T_1993;
  wire [15:0] _T_1994;
  wire [1:0] _T_1995;
  wire [1:0] _T_1996;
  wire [3:0] _T_1997;
  wire [1:0] _T_1998;
  wire [1:0] _T_1999;
  wire [3:0] _T_2000;
  wire [7:0] _T_2001;
  wire [1:0] _T_2002;
  wire [1:0] _T_2003;
  wire [3:0] _T_2004;
  wire [1:0] _T_2005;
  wire [1:0] _T_2006;
  wire [3:0] _T_2007;
  wire [7:0] _T_2008;
  wire [15:0] _T_2009;
  wire [31:0] _T_2010;
  wire [1:0] _T_2011;
  wire [1:0] _T_2012;
  wire [3:0] _T_2013;
  wire [1:0] _T_2014;
  wire [1:0] _T_2015;
  wire [3:0] _T_2016;
  wire [7:0] _T_2017;
  wire [1:0] _T_2018;
  wire [1:0] _T_2019;
  wire [3:0] _T_2020;
  wire [1:0] _T_2021;
  wire [1:0] _T_2022;
  wire [3:0] _T_2023;
  wire [7:0] _T_2024;
  wire [15:0] _T_2025;
  wire [1:0] _T_2026;
  wire [1:0] _T_2027;
  wire [3:0] _T_2028;
  wire [1:0] _T_2029;
  wire [1:0] _T_2030;
  wire [3:0] _T_2031;
  wire [7:0] _T_2032;
  wire [1:0] _T_2033;
  wire [1:0] _T_2034;
  wire [3:0] _T_2035;
  wire [1:0] _T_2036;
  wire [1:0] _T_2037;
  wire [3:0] _T_2038;
  wire [7:0] _T_2039;
  wire [15:0] _T_2040;
  wire [31:0] _T_2041;
  wire [63:0] _T_2042;
  wire [1:0] _T_2043;
  wire [1:0] _T_2044;
  wire [3:0] _T_2045;
  wire [1:0] _T_2046;
  wire [1:0] _T_2047;
  wire [3:0] _T_2048;
  wire [7:0] _T_2049;
  wire [1:0] _T_2050;
  wire [1:0] _T_2051;
  wire [3:0] _T_2052;
  wire [1:0] _T_2053;
  wire [1:0] _T_2054;
  wire [3:0] _T_2055;
  wire [7:0] _T_2056;
  wire [15:0] _T_2057;
  wire [1:0] _T_2058;
  wire [1:0] _T_2059;
  wire [3:0] _T_2060;
  wire [1:0] _T_2061;
  wire [1:0] _T_2062;
  wire [3:0] _T_2063;
  wire [7:0] _T_2064;
  wire [1:0] _T_2065;
  wire [1:0] _T_2066;
  wire [3:0] _T_2067;
  wire [1:0] _T_2068;
  wire [1:0] _T_2069;
  wire [3:0] _T_2070;
  wire [7:0] _T_2071;
  wire [15:0] _T_2072;
  wire [31:0] _T_2073;
  wire [1:0] _T_2074;
  wire [1:0] _T_2075;
  wire [3:0] _T_2076;
  wire [1:0] _T_2077;
  wire [1:0] _T_2078;
  wire [3:0] _T_2079;
  wire [7:0] _T_2080;
  wire [1:0] _T_2081;
  wire [1:0] _T_2082;
  wire [3:0] _T_2083;
  wire [1:0] _T_2084;
  wire [1:0] _T_2085;
  wire [3:0] _T_2086;
  wire [7:0] _T_2087;
  wire [15:0] _T_2088;
  wire [1:0] _T_2089;
  wire [1:0] _T_2090;
  wire [3:0] _T_2091;
  wire [1:0] _T_2092;
  wire [1:0] _T_2093;
  wire [3:0] _T_2094;
  wire [7:0] _T_2095;
  wire [1:0] _T_2096;
  wire [1:0] _T_2097;
  wire [3:0] _T_2098;
  wire [1:0] _T_2099;
  wire [1:0] _T_2100;
  wire [3:0] _T_2101;
  wire [7:0] _T_2102;
  wire [15:0] _T_2103;
  wire [31:0] _T_2104;
  wire [63:0] _T_2105;
  wire [127:0] _T_2106;
  wire [255:0] _T_2107;
  wire [511:0] _T_2108;
  wire  _T_2113;
  wire  _T_2114;
  wire [9:0] _GEN_1538;
  assign io_inputMemConsumed = _T_1056;
  assign io_outputMemBlock = _T_2108;
  assign io_outputMemBlockValid = _T_1597;
  assign io_outputBits = outputBits;
  assign io_outputFinished = _T_2114;
  assign _T_540 = io_inputMemBlock[0];
  assign _T_541 = io_inputMemBlock[1];
  assign _T_542 = io_inputMemBlock[2];
  assign _T_543 = io_inputMemBlock[3];
  assign _T_544 = io_inputMemBlock[4];
  assign _T_545 = io_inputMemBlock[5];
  assign _T_546 = io_inputMemBlock[6];
  assign _T_547 = io_inputMemBlock[7];
  assign _T_548 = io_inputMemBlock[8];
  assign _T_549 = io_inputMemBlock[9];
  assign _T_550 = io_inputMemBlock[10];
  assign _T_551 = io_inputMemBlock[11];
  assign _T_552 = io_inputMemBlock[12];
  assign _T_553 = io_inputMemBlock[13];
  assign _T_554 = io_inputMemBlock[14];
  assign _T_555 = io_inputMemBlock[15];
  assign _T_556 = io_inputMemBlock[16];
  assign _T_557 = io_inputMemBlock[17];
  assign _T_558 = io_inputMemBlock[18];
  assign _T_559 = io_inputMemBlock[19];
  assign _T_560 = io_inputMemBlock[20];
  assign _T_561 = io_inputMemBlock[21];
  assign _T_562 = io_inputMemBlock[22];
  assign _T_563 = io_inputMemBlock[23];
  assign _T_564 = io_inputMemBlock[24];
  assign _T_565 = io_inputMemBlock[25];
  assign _T_566 = io_inputMemBlock[26];
  assign _T_567 = io_inputMemBlock[27];
  assign _T_568 = io_inputMemBlock[28];
  assign _T_569 = io_inputMemBlock[29];
  assign _T_570 = io_inputMemBlock[30];
  assign _T_571 = io_inputMemBlock[31];
  assign _T_572 = io_inputMemBlock[32];
  assign _T_573 = io_inputMemBlock[33];
  assign _T_574 = io_inputMemBlock[34];
  assign _T_575 = io_inputMemBlock[35];
  assign _T_576 = io_inputMemBlock[36];
  assign _T_577 = io_inputMemBlock[37];
  assign _T_578 = io_inputMemBlock[38];
  assign _T_579 = io_inputMemBlock[39];
  assign _T_580 = io_inputMemBlock[40];
  assign _T_581 = io_inputMemBlock[41];
  assign _T_582 = io_inputMemBlock[42];
  assign _T_583 = io_inputMemBlock[43];
  assign _T_584 = io_inputMemBlock[44];
  assign _T_585 = io_inputMemBlock[45];
  assign _T_586 = io_inputMemBlock[46];
  assign _T_587 = io_inputMemBlock[47];
  assign _T_588 = io_inputMemBlock[48];
  assign _T_589 = io_inputMemBlock[49];
  assign _T_590 = io_inputMemBlock[50];
  assign _T_591 = io_inputMemBlock[51];
  assign _T_592 = io_inputMemBlock[52];
  assign _T_593 = io_inputMemBlock[53];
  assign _T_594 = io_inputMemBlock[54];
  assign _T_595 = io_inputMemBlock[55];
  assign _T_596 = io_inputMemBlock[56];
  assign _T_597 = io_inputMemBlock[57];
  assign _T_598 = io_inputMemBlock[58];
  assign _T_599 = io_inputMemBlock[59];
  assign _T_600 = io_inputMemBlock[60];
  assign _T_601 = io_inputMemBlock[61];
  assign _T_602 = io_inputMemBlock[62];
  assign _T_603 = io_inputMemBlock[63];
  assign _T_604 = io_inputMemBlock[64];
  assign _T_605 = io_inputMemBlock[65];
  assign _T_606 = io_inputMemBlock[66];
  assign _T_607 = io_inputMemBlock[67];
  assign _T_608 = io_inputMemBlock[68];
  assign _T_609 = io_inputMemBlock[69];
  assign _T_610 = io_inputMemBlock[70];
  assign _T_611 = io_inputMemBlock[71];
  assign _T_612 = io_inputMemBlock[72];
  assign _T_613 = io_inputMemBlock[73];
  assign _T_614 = io_inputMemBlock[74];
  assign _T_615 = io_inputMemBlock[75];
  assign _T_616 = io_inputMemBlock[76];
  assign _T_617 = io_inputMemBlock[77];
  assign _T_618 = io_inputMemBlock[78];
  assign _T_619 = io_inputMemBlock[79];
  assign _T_620 = io_inputMemBlock[80];
  assign _T_621 = io_inputMemBlock[81];
  assign _T_622 = io_inputMemBlock[82];
  assign _T_623 = io_inputMemBlock[83];
  assign _T_624 = io_inputMemBlock[84];
  assign _T_625 = io_inputMemBlock[85];
  assign _T_626 = io_inputMemBlock[86];
  assign _T_627 = io_inputMemBlock[87];
  assign _T_628 = io_inputMemBlock[88];
  assign _T_629 = io_inputMemBlock[89];
  assign _T_630 = io_inputMemBlock[90];
  assign _T_631 = io_inputMemBlock[91];
  assign _T_632 = io_inputMemBlock[92];
  assign _T_633 = io_inputMemBlock[93];
  assign _T_634 = io_inputMemBlock[94];
  assign _T_635 = io_inputMemBlock[95];
  assign _T_636 = io_inputMemBlock[96];
  assign _T_637 = io_inputMemBlock[97];
  assign _T_638 = io_inputMemBlock[98];
  assign _T_639 = io_inputMemBlock[99];
  assign _T_640 = io_inputMemBlock[100];
  assign _T_641 = io_inputMemBlock[101];
  assign _T_642 = io_inputMemBlock[102];
  assign _T_643 = io_inputMemBlock[103];
  assign _T_644 = io_inputMemBlock[104];
  assign _T_645 = io_inputMemBlock[105];
  assign _T_646 = io_inputMemBlock[106];
  assign _T_647 = io_inputMemBlock[107];
  assign _T_648 = io_inputMemBlock[108];
  assign _T_649 = io_inputMemBlock[109];
  assign _T_650 = io_inputMemBlock[110];
  assign _T_651 = io_inputMemBlock[111];
  assign _T_652 = io_inputMemBlock[112];
  assign _T_653 = io_inputMemBlock[113];
  assign _T_654 = io_inputMemBlock[114];
  assign _T_655 = io_inputMemBlock[115];
  assign _T_656 = io_inputMemBlock[116];
  assign _T_657 = io_inputMemBlock[117];
  assign _T_658 = io_inputMemBlock[118];
  assign _T_659 = io_inputMemBlock[119];
  assign _T_660 = io_inputMemBlock[120];
  assign _T_661 = io_inputMemBlock[121];
  assign _T_662 = io_inputMemBlock[122];
  assign _T_663 = io_inputMemBlock[123];
  assign _T_664 = io_inputMemBlock[124];
  assign _T_665 = io_inputMemBlock[125];
  assign _T_666 = io_inputMemBlock[126];
  assign _T_667 = io_inputMemBlock[127];
  assign _T_668 = io_inputMemBlock[128];
  assign _T_669 = io_inputMemBlock[129];
  assign _T_670 = io_inputMemBlock[130];
  assign _T_671 = io_inputMemBlock[131];
  assign _T_672 = io_inputMemBlock[132];
  assign _T_673 = io_inputMemBlock[133];
  assign _T_674 = io_inputMemBlock[134];
  assign _T_675 = io_inputMemBlock[135];
  assign _T_676 = io_inputMemBlock[136];
  assign _T_677 = io_inputMemBlock[137];
  assign _T_678 = io_inputMemBlock[138];
  assign _T_679 = io_inputMemBlock[139];
  assign _T_680 = io_inputMemBlock[140];
  assign _T_681 = io_inputMemBlock[141];
  assign _T_682 = io_inputMemBlock[142];
  assign _T_683 = io_inputMemBlock[143];
  assign _T_684 = io_inputMemBlock[144];
  assign _T_685 = io_inputMemBlock[145];
  assign _T_686 = io_inputMemBlock[146];
  assign _T_687 = io_inputMemBlock[147];
  assign _T_688 = io_inputMemBlock[148];
  assign _T_689 = io_inputMemBlock[149];
  assign _T_690 = io_inputMemBlock[150];
  assign _T_691 = io_inputMemBlock[151];
  assign _T_692 = io_inputMemBlock[152];
  assign _T_693 = io_inputMemBlock[153];
  assign _T_694 = io_inputMemBlock[154];
  assign _T_695 = io_inputMemBlock[155];
  assign _T_696 = io_inputMemBlock[156];
  assign _T_697 = io_inputMemBlock[157];
  assign _T_698 = io_inputMemBlock[158];
  assign _T_699 = io_inputMemBlock[159];
  assign _T_700 = io_inputMemBlock[160];
  assign _T_701 = io_inputMemBlock[161];
  assign _T_702 = io_inputMemBlock[162];
  assign _T_703 = io_inputMemBlock[163];
  assign _T_704 = io_inputMemBlock[164];
  assign _T_705 = io_inputMemBlock[165];
  assign _T_706 = io_inputMemBlock[166];
  assign _T_707 = io_inputMemBlock[167];
  assign _T_708 = io_inputMemBlock[168];
  assign _T_709 = io_inputMemBlock[169];
  assign _T_710 = io_inputMemBlock[170];
  assign _T_711 = io_inputMemBlock[171];
  assign _T_712 = io_inputMemBlock[172];
  assign _T_713 = io_inputMemBlock[173];
  assign _T_714 = io_inputMemBlock[174];
  assign _T_715 = io_inputMemBlock[175];
  assign _T_716 = io_inputMemBlock[176];
  assign _T_717 = io_inputMemBlock[177];
  assign _T_718 = io_inputMemBlock[178];
  assign _T_719 = io_inputMemBlock[179];
  assign _T_720 = io_inputMemBlock[180];
  assign _T_721 = io_inputMemBlock[181];
  assign _T_722 = io_inputMemBlock[182];
  assign _T_723 = io_inputMemBlock[183];
  assign _T_724 = io_inputMemBlock[184];
  assign _T_725 = io_inputMemBlock[185];
  assign _T_726 = io_inputMemBlock[186];
  assign _T_727 = io_inputMemBlock[187];
  assign _T_728 = io_inputMemBlock[188];
  assign _T_729 = io_inputMemBlock[189];
  assign _T_730 = io_inputMemBlock[190];
  assign _T_731 = io_inputMemBlock[191];
  assign _T_732 = io_inputMemBlock[192];
  assign _T_733 = io_inputMemBlock[193];
  assign _T_734 = io_inputMemBlock[194];
  assign _T_735 = io_inputMemBlock[195];
  assign _T_736 = io_inputMemBlock[196];
  assign _T_737 = io_inputMemBlock[197];
  assign _T_738 = io_inputMemBlock[198];
  assign _T_739 = io_inputMemBlock[199];
  assign _T_740 = io_inputMemBlock[200];
  assign _T_741 = io_inputMemBlock[201];
  assign _T_742 = io_inputMemBlock[202];
  assign _T_743 = io_inputMemBlock[203];
  assign _T_744 = io_inputMemBlock[204];
  assign _T_745 = io_inputMemBlock[205];
  assign _T_746 = io_inputMemBlock[206];
  assign _T_747 = io_inputMemBlock[207];
  assign _T_748 = io_inputMemBlock[208];
  assign _T_749 = io_inputMemBlock[209];
  assign _T_750 = io_inputMemBlock[210];
  assign _T_751 = io_inputMemBlock[211];
  assign _T_752 = io_inputMemBlock[212];
  assign _T_753 = io_inputMemBlock[213];
  assign _T_754 = io_inputMemBlock[214];
  assign _T_755 = io_inputMemBlock[215];
  assign _T_756 = io_inputMemBlock[216];
  assign _T_757 = io_inputMemBlock[217];
  assign _T_758 = io_inputMemBlock[218];
  assign _T_759 = io_inputMemBlock[219];
  assign _T_760 = io_inputMemBlock[220];
  assign _T_761 = io_inputMemBlock[221];
  assign _T_762 = io_inputMemBlock[222];
  assign _T_763 = io_inputMemBlock[223];
  assign _T_764 = io_inputMemBlock[224];
  assign _T_765 = io_inputMemBlock[225];
  assign _T_766 = io_inputMemBlock[226];
  assign _T_767 = io_inputMemBlock[227];
  assign _T_768 = io_inputMemBlock[228];
  assign _T_769 = io_inputMemBlock[229];
  assign _T_770 = io_inputMemBlock[230];
  assign _T_771 = io_inputMemBlock[231];
  assign _T_772 = io_inputMemBlock[232];
  assign _T_773 = io_inputMemBlock[233];
  assign _T_774 = io_inputMemBlock[234];
  assign _T_775 = io_inputMemBlock[235];
  assign _T_776 = io_inputMemBlock[236];
  assign _T_777 = io_inputMemBlock[237];
  assign _T_778 = io_inputMemBlock[238];
  assign _T_779 = io_inputMemBlock[239];
  assign _T_780 = io_inputMemBlock[240];
  assign _T_781 = io_inputMemBlock[241];
  assign _T_782 = io_inputMemBlock[242];
  assign _T_783 = io_inputMemBlock[243];
  assign _T_784 = io_inputMemBlock[244];
  assign _T_785 = io_inputMemBlock[245];
  assign _T_786 = io_inputMemBlock[246];
  assign _T_787 = io_inputMemBlock[247];
  assign _T_788 = io_inputMemBlock[248];
  assign _T_789 = io_inputMemBlock[249];
  assign _T_790 = io_inputMemBlock[250];
  assign _T_791 = io_inputMemBlock[251];
  assign _T_792 = io_inputMemBlock[252];
  assign _T_793 = io_inputMemBlock[253];
  assign _T_794 = io_inputMemBlock[254];
  assign _T_795 = io_inputMemBlock[255];
  assign _T_796 = io_inputMemBlock[256];
  assign _T_797 = io_inputMemBlock[257];
  assign _T_798 = io_inputMemBlock[258];
  assign _T_799 = io_inputMemBlock[259];
  assign _T_800 = io_inputMemBlock[260];
  assign _T_801 = io_inputMemBlock[261];
  assign _T_802 = io_inputMemBlock[262];
  assign _T_803 = io_inputMemBlock[263];
  assign _T_804 = io_inputMemBlock[264];
  assign _T_805 = io_inputMemBlock[265];
  assign _T_806 = io_inputMemBlock[266];
  assign _T_807 = io_inputMemBlock[267];
  assign _T_808 = io_inputMemBlock[268];
  assign _T_809 = io_inputMemBlock[269];
  assign _T_810 = io_inputMemBlock[270];
  assign _T_811 = io_inputMemBlock[271];
  assign _T_812 = io_inputMemBlock[272];
  assign _T_813 = io_inputMemBlock[273];
  assign _T_814 = io_inputMemBlock[274];
  assign _T_815 = io_inputMemBlock[275];
  assign _T_816 = io_inputMemBlock[276];
  assign _T_817 = io_inputMemBlock[277];
  assign _T_818 = io_inputMemBlock[278];
  assign _T_819 = io_inputMemBlock[279];
  assign _T_820 = io_inputMemBlock[280];
  assign _T_821 = io_inputMemBlock[281];
  assign _T_822 = io_inputMemBlock[282];
  assign _T_823 = io_inputMemBlock[283];
  assign _T_824 = io_inputMemBlock[284];
  assign _T_825 = io_inputMemBlock[285];
  assign _T_826 = io_inputMemBlock[286];
  assign _T_827 = io_inputMemBlock[287];
  assign _T_828 = io_inputMemBlock[288];
  assign _T_829 = io_inputMemBlock[289];
  assign _T_830 = io_inputMemBlock[290];
  assign _T_831 = io_inputMemBlock[291];
  assign _T_832 = io_inputMemBlock[292];
  assign _T_833 = io_inputMemBlock[293];
  assign _T_834 = io_inputMemBlock[294];
  assign _T_835 = io_inputMemBlock[295];
  assign _T_836 = io_inputMemBlock[296];
  assign _T_837 = io_inputMemBlock[297];
  assign _T_838 = io_inputMemBlock[298];
  assign _T_839 = io_inputMemBlock[299];
  assign _T_840 = io_inputMemBlock[300];
  assign _T_841 = io_inputMemBlock[301];
  assign _T_842 = io_inputMemBlock[302];
  assign _T_843 = io_inputMemBlock[303];
  assign _T_844 = io_inputMemBlock[304];
  assign _T_845 = io_inputMemBlock[305];
  assign _T_846 = io_inputMemBlock[306];
  assign _T_847 = io_inputMemBlock[307];
  assign _T_848 = io_inputMemBlock[308];
  assign _T_849 = io_inputMemBlock[309];
  assign _T_850 = io_inputMemBlock[310];
  assign _T_851 = io_inputMemBlock[311];
  assign _T_852 = io_inputMemBlock[312];
  assign _T_853 = io_inputMemBlock[313];
  assign _T_854 = io_inputMemBlock[314];
  assign _T_855 = io_inputMemBlock[315];
  assign _T_856 = io_inputMemBlock[316];
  assign _T_857 = io_inputMemBlock[317];
  assign _T_858 = io_inputMemBlock[318];
  assign _T_859 = io_inputMemBlock[319];
  assign _T_860 = io_inputMemBlock[320];
  assign _T_861 = io_inputMemBlock[321];
  assign _T_862 = io_inputMemBlock[322];
  assign _T_863 = io_inputMemBlock[323];
  assign _T_864 = io_inputMemBlock[324];
  assign _T_865 = io_inputMemBlock[325];
  assign _T_866 = io_inputMemBlock[326];
  assign _T_867 = io_inputMemBlock[327];
  assign _T_868 = io_inputMemBlock[328];
  assign _T_869 = io_inputMemBlock[329];
  assign _T_870 = io_inputMemBlock[330];
  assign _T_871 = io_inputMemBlock[331];
  assign _T_872 = io_inputMemBlock[332];
  assign _T_873 = io_inputMemBlock[333];
  assign _T_874 = io_inputMemBlock[334];
  assign _T_875 = io_inputMemBlock[335];
  assign _T_876 = io_inputMemBlock[336];
  assign _T_877 = io_inputMemBlock[337];
  assign _T_878 = io_inputMemBlock[338];
  assign _T_879 = io_inputMemBlock[339];
  assign _T_880 = io_inputMemBlock[340];
  assign _T_881 = io_inputMemBlock[341];
  assign _T_882 = io_inputMemBlock[342];
  assign _T_883 = io_inputMemBlock[343];
  assign _T_884 = io_inputMemBlock[344];
  assign _T_885 = io_inputMemBlock[345];
  assign _T_886 = io_inputMemBlock[346];
  assign _T_887 = io_inputMemBlock[347];
  assign _T_888 = io_inputMemBlock[348];
  assign _T_889 = io_inputMemBlock[349];
  assign _T_890 = io_inputMemBlock[350];
  assign _T_891 = io_inputMemBlock[351];
  assign _T_892 = io_inputMemBlock[352];
  assign _T_893 = io_inputMemBlock[353];
  assign _T_894 = io_inputMemBlock[354];
  assign _T_895 = io_inputMemBlock[355];
  assign _T_896 = io_inputMemBlock[356];
  assign _T_897 = io_inputMemBlock[357];
  assign _T_898 = io_inputMemBlock[358];
  assign _T_899 = io_inputMemBlock[359];
  assign _T_900 = io_inputMemBlock[360];
  assign _T_901 = io_inputMemBlock[361];
  assign _T_902 = io_inputMemBlock[362];
  assign _T_903 = io_inputMemBlock[363];
  assign _T_904 = io_inputMemBlock[364];
  assign _T_905 = io_inputMemBlock[365];
  assign _T_906 = io_inputMemBlock[366];
  assign _T_907 = io_inputMemBlock[367];
  assign _T_908 = io_inputMemBlock[368];
  assign _T_909 = io_inputMemBlock[369];
  assign _T_910 = io_inputMemBlock[370];
  assign _T_911 = io_inputMemBlock[371];
  assign _T_912 = io_inputMemBlock[372];
  assign _T_913 = io_inputMemBlock[373];
  assign _T_914 = io_inputMemBlock[374];
  assign _T_915 = io_inputMemBlock[375];
  assign _T_916 = io_inputMemBlock[376];
  assign _T_917 = io_inputMemBlock[377];
  assign _T_918 = io_inputMemBlock[378];
  assign _T_919 = io_inputMemBlock[379];
  assign _T_920 = io_inputMemBlock[380];
  assign _T_921 = io_inputMemBlock[381];
  assign _T_922 = io_inputMemBlock[382];
  assign _T_923 = io_inputMemBlock[383];
  assign _T_924 = io_inputMemBlock[384];
  assign _T_925 = io_inputMemBlock[385];
  assign _T_926 = io_inputMemBlock[386];
  assign _T_927 = io_inputMemBlock[387];
  assign _T_928 = io_inputMemBlock[388];
  assign _T_929 = io_inputMemBlock[389];
  assign _T_930 = io_inputMemBlock[390];
  assign _T_931 = io_inputMemBlock[391];
  assign _T_932 = io_inputMemBlock[392];
  assign _T_933 = io_inputMemBlock[393];
  assign _T_934 = io_inputMemBlock[394];
  assign _T_935 = io_inputMemBlock[395];
  assign _T_936 = io_inputMemBlock[396];
  assign _T_937 = io_inputMemBlock[397];
  assign _T_938 = io_inputMemBlock[398];
  assign _T_939 = io_inputMemBlock[399];
  assign _T_940 = io_inputMemBlock[400];
  assign _T_941 = io_inputMemBlock[401];
  assign _T_942 = io_inputMemBlock[402];
  assign _T_943 = io_inputMemBlock[403];
  assign _T_944 = io_inputMemBlock[404];
  assign _T_945 = io_inputMemBlock[405];
  assign _T_946 = io_inputMemBlock[406];
  assign _T_947 = io_inputMemBlock[407];
  assign _T_948 = io_inputMemBlock[408];
  assign _T_949 = io_inputMemBlock[409];
  assign _T_950 = io_inputMemBlock[410];
  assign _T_951 = io_inputMemBlock[411];
  assign _T_952 = io_inputMemBlock[412];
  assign _T_953 = io_inputMemBlock[413];
  assign _T_954 = io_inputMemBlock[414];
  assign _T_955 = io_inputMemBlock[415];
  assign _T_956 = io_inputMemBlock[416];
  assign _T_957 = io_inputMemBlock[417];
  assign _T_958 = io_inputMemBlock[418];
  assign _T_959 = io_inputMemBlock[419];
  assign _T_960 = io_inputMemBlock[420];
  assign _T_961 = io_inputMemBlock[421];
  assign _T_962 = io_inputMemBlock[422];
  assign _T_963 = io_inputMemBlock[423];
  assign _T_964 = io_inputMemBlock[424];
  assign _T_965 = io_inputMemBlock[425];
  assign _T_966 = io_inputMemBlock[426];
  assign _T_967 = io_inputMemBlock[427];
  assign _T_968 = io_inputMemBlock[428];
  assign _T_969 = io_inputMemBlock[429];
  assign _T_970 = io_inputMemBlock[430];
  assign _T_971 = io_inputMemBlock[431];
  assign _T_972 = io_inputMemBlock[432];
  assign _T_973 = io_inputMemBlock[433];
  assign _T_974 = io_inputMemBlock[434];
  assign _T_975 = io_inputMemBlock[435];
  assign _T_976 = io_inputMemBlock[436];
  assign _T_977 = io_inputMemBlock[437];
  assign _T_978 = io_inputMemBlock[438];
  assign _T_979 = io_inputMemBlock[439];
  assign _T_980 = io_inputMemBlock[440];
  assign _T_981 = io_inputMemBlock[441];
  assign _T_982 = io_inputMemBlock[442];
  assign _T_983 = io_inputMemBlock[443];
  assign _T_984 = io_inputMemBlock[444];
  assign _T_985 = io_inputMemBlock[445];
  assign _T_986 = io_inputMemBlock[446];
  assign _T_987 = io_inputMemBlock[447];
  assign _T_988 = io_inputMemBlock[448];
  assign _T_989 = io_inputMemBlock[449];
  assign _T_990 = io_inputMemBlock[450];
  assign _T_991 = io_inputMemBlock[451];
  assign _T_992 = io_inputMemBlock[452];
  assign _T_993 = io_inputMemBlock[453];
  assign _T_994 = io_inputMemBlock[454];
  assign _T_995 = io_inputMemBlock[455];
  assign _T_996 = io_inputMemBlock[456];
  assign _T_997 = io_inputMemBlock[457];
  assign _T_998 = io_inputMemBlock[458];
  assign _T_999 = io_inputMemBlock[459];
  assign _T_1000 = io_inputMemBlock[460];
  assign _T_1001 = io_inputMemBlock[461];
  assign _T_1002 = io_inputMemBlock[462];
  assign _T_1003 = io_inputMemBlock[463];
  assign _T_1004 = io_inputMemBlock[464];
  assign _T_1005 = io_inputMemBlock[465];
  assign _T_1006 = io_inputMemBlock[466];
  assign _T_1007 = io_inputMemBlock[467];
  assign _T_1008 = io_inputMemBlock[468];
  assign _T_1009 = io_inputMemBlock[469];
  assign _T_1010 = io_inputMemBlock[470];
  assign _T_1011 = io_inputMemBlock[471];
  assign _T_1012 = io_inputMemBlock[472];
  assign _T_1013 = io_inputMemBlock[473];
  assign _T_1014 = io_inputMemBlock[474];
  assign _T_1015 = io_inputMemBlock[475];
  assign _T_1016 = io_inputMemBlock[476];
  assign _T_1017 = io_inputMemBlock[477];
  assign _T_1018 = io_inputMemBlock[478];
  assign _T_1019 = io_inputMemBlock[479];
  assign _T_1020 = io_inputMemBlock[480];
  assign _T_1021 = io_inputMemBlock[481];
  assign _T_1022 = io_inputMemBlock[482];
  assign _T_1023 = io_inputMemBlock[483];
  assign _T_1024 = io_inputMemBlock[484];
  assign _T_1025 = io_inputMemBlock[485];
  assign _T_1026 = io_inputMemBlock[486];
  assign _T_1027 = io_inputMemBlock[487];
  assign _T_1028 = io_inputMemBlock[488];
  assign _T_1029 = io_inputMemBlock[489];
  assign _T_1030 = io_inputMemBlock[490];
  assign _T_1031 = io_inputMemBlock[491];
  assign _T_1032 = io_inputMemBlock[492];
  assign _T_1033 = io_inputMemBlock[493];
  assign _T_1034 = io_inputMemBlock[494];
  assign _T_1035 = io_inputMemBlock[495];
  assign _T_1036 = io_inputMemBlock[496];
  assign _T_1037 = io_inputMemBlock[497];
  assign _T_1038 = io_inputMemBlock[498];
  assign _T_1039 = io_inputMemBlock[499];
  assign _T_1040 = io_inputMemBlock[500];
  assign _T_1041 = io_inputMemBlock[501];
  assign _T_1042 = io_inputMemBlock[502];
  assign _T_1043 = io_inputMemBlock[503];
  assign _T_1044 = io_inputMemBlock[504];
  assign _T_1045 = io_inputMemBlock[505];
  assign _T_1046 = io_inputMemBlock[506];
  assign _T_1047 = io_inputMemBlock[507];
  assign _T_1048 = io_inputMemBlock[508];
  assign _T_1049 = io_inputMemBlock[509];
  assign _T_1050 = io_inputMemBlock[510];
  assign _T_1051 = io_inputMemBlock[511];
  assign _GEN_0 = io_inputMemBlockValid ? io_inputBits : inputBitsRemaining;
  assign _GEN_1 = io_inputMemBlockValid ? _T_540 : inputMemBlock_0;
  assign _GEN_2 = io_inputMemBlockValid ? _T_541 : inputMemBlock_1;
  assign _GEN_3 = io_inputMemBlockValid ? _T_542 : inputMemBlock_2;
  assign _GEN_4 = io_inputMemBlockValid ? _T_543 : inputMemBlock_3;
  assign _GEN_5 = io_inputMemBlockValid ? _T_544 : inputMemBlock_4;
  assign _GEN_6 = io_inputMemBlockValid ? _T_545 : inputMemBlock_5;
  assign _GEN_7 = io_inputMemBlockValid ? _T_546 : inputMemBlock_6;
  assign _GEN_8 = io_inputMemBlockValid ? _T_547 : inputMemBlock_7;
  assign _GEN_9 = io_inputMemBlockValid ? _T_548 : inputMemBlock_8;
  assign _GEN_10 = io_inputMemBlockValid ? _T_549 : inputMemBlock_9;
  assign _GEN_11 = io_inputMemBlockValid ? _T_550 : inputMemBlock_10;
  assign _GEN_12 = io_inputMemBlockValid ? _T_551 : inputMemBlock_11;
  assign _GEN_13 = io_inputMemBlockValid ? _T_552 : inputMemBlock_12;
  assign _GEN_14 = io_inputMemBlockValid ? _T_553 : inputMemBlock_13;
  assign _GEN_15 = io_inputMemBlockValid ? _T_554 : inputMemBlock_14;
  assign _GEN_16 = io_inputMemBlockValid ? _T_555 : inputMemBlock_15;
  assign _GEN_17 = io_inputMemBlockValid ? _T_556 : inputMemBlock_16;
  assign _GEN_18 = io_inputMemBlockValid ? _T_557 : inputMemBlock_17;
  assign _GEN_19 = io_inputMemBlockValid ? _T_558 : inputMemBlock_18;
  assign _GEN_20 = io_inputMemBlockValid ? _T_559 : inputMemBlock_19;
  assign _GEN_21 = io_inputMemBlockValid ? _T_560 : inputMemBlock_20;
  assign _GEN_22 = io_inputMemBlockValid ? _T_561 : inputMemBlock_21;
  assign _GEN_23 = io_inputMemBlockValid ? _T_562 : inputMemBlock_22;
  assign _GEN_24 = io_inputMemBlockValid ? _T_563 : inputMemBlock_23;
  assign _GEN_25 = io_inputMemBlockValid ? _T_564 : inputMemBlock_24;
  assign _GEN_26 = io_inputMemBlockValid ? _T_565 : inputMemBlock_25;
  assign _GEN_27 = io_inputMemBlockValid ? _T_566 : inputMemBlock_26;
  assign _GEN_28 = io_inputMemBlockValid ? _T_567 : inputMemBlock_27;
  assign _GEN_29 = io_inputMemBlockValid ? _T_568 : inputMemBlock_28;
  assign _GEN_30 = io_inputMemBlockValid ? _T_569 : inputMemBlock_29;
  assign _GEN_31 = io_inputMemBlockValid ? _T_570 : inputMemBlock_30;
  assign _GEN_32 = io_inputMemBlockValid ? _T_571 : inputMemBlock_31;
  assign _GEN_33 = io_inputMemBlockValid ? _T_572 : inputMemBlock_32;
  assign _GEN_34 = io_inputMemBlockValid ? _T_573 : inputMemBlock_33;
  assign _GEN_35 = io_inputMemBlockValid ? _T_574 : inputMemBlock_34;
  assign _GEN_36 = io_inputMemBlockValid ? _T_575 : inputMemBlock_35;
  assign _GEN_37 = io_inputMemBlockValid ? _T_576 : inputMemBlock_36;
  assign _GEN_38 = io_inputMemBlockValid ? _T_577 : inputMemBlock_37;
  assign _GEN_39 = io_inputMemBlockValid ? _T_578 : inputMemBlock_38;
  assign _GEN_40 = io_inputMemBlockValid ? _T_579 : inputMemBlock_39;
  assign _GEN_41 = io_inputMemBlockValid ? _T_580 : inputMemBlock_40;
  assign _GEN_42 = io_inputMemBlockValid ? _T_581 : inputMemBlock_41;
  assign _GEN_43 = io_inputMemBlockValid ? _T_582 : inputMemBlock_42;
  assign _GEN_44 = io_inputMemBlockValid ? _T_583 : inputMemBlock_43;
  assign _GEN_45 = io_inputMemBlockValid ? _T_584 : inputMemBlock_44;
  assign _GEN_46 = io_inputMemBlockValid ? _T_585 : inputMemBlock_45;
  assign _GEN_47 = io_inputMemBlockValid ? _T_586 : inputMemBlock_46;
  assign _GEN_48 = io_inputMemBlockValid ? _T_587 : inputMemBlock_47;
  assign _GEN_49 = io_inputMemBlockValid ? _T_588 : inputMemBlock_48;
  assign _GEN_50 = io_inputMemBlockValid ? _T_589 : inputMemBlock_49;
  assign _GEN_51 = io_inputMemBlockValid ? _T_590 : inputMemBlock_50;
  assign _GEN_52 = io_inputMemBlockValid ? _T_591 : inputMemBlock_51;
  assign _GEN_53 = io_inputMemBlockValid ? _T_592 : inputMemBlock_52;
  assign _GEN_54 = io_inputMemBlockValid ? _T_593 : inputMemBlock_53;
  assign _GEN_55 = io_inputMemBlockValid ? _T_594 : inputMemBlock_54;
  assign _GEN_56 = io_inputMemBlockValid ? _T_595 : inputMemBlock_55;
  assign _GEN_57 = io_inputMemBlockValid ? _T_596 : inputMemBlock_56;
  assign _GEN_58 = io_inputMemBlockValid ? _T_597 : inputMemBlock_57;
  assign _GEN_59 = io_inputMemBlockValid ? _T_598 : inputMemBlock_58;
  assign _GEN_60 = io_inputMemBlockValid ? _T_599 : inputMemBlock_59;
  assign _GEN_61 = io_inputMemBlockValid ? _T_600 : inputMemBlock_60;
  assign _GEN_62 = io_inputMemBlockValid ? _T_601 : inputMemBlock_61;
  assign _GEN_63 = io_inputMemBlockValid ? _T_602 : inputMemBlock_62;
  assign _GEN_64 = io_inputMemBlockValid ? _T_603 : inputMemBlock_63;
  assign _GEN_65 = io_inputMemBlockValid ? _T_604 : inputMemBlock_64;
  assign _GEN_66 = io_inputMemBlockValid ? _T_605 : inputMemBlock_65;
  assign _GEN_67 = io_inputMemBlockValid ? _T_606 : inputMemBlock_66;
  assign _GEN_68 = io_inputMemBlockValid ? _T_607 : inputMemBlock_67;
  assign _GEN_69 = io_inputMemBlockValid ? _T_608 : inputMemBlock_68;
  assign _GEN_70 = io_inputMemBlockValid ? _T_609 : inputMemBlock_69;
  assign _GEN_71 = io_inputMemBlockValid ? _T_610 : inputMemBlock_70;
  assign _GEN_72 = io_inputMemBlockValid ? _T_611 : inputMemBlock_71;
  assign _GEN_73 = io_inputMemBlockValid ? _T_612 : inputMemBlock_72;
  assign _GEN_74 = io_inputMemBlockValid ? _T_613 : inputMemBlock_73;
  assign _GEN_75 = io_inputMemBlockValid ? _T_614 : inputMemBlock_74;
  assign _GEN_76 = io_inputMemBlockValid ? _T_615 : inputMemBlock_75;
  assign _GEN_77 = io_inputMemBlockValid ? _T_616 : inputMemBlock_76;
  assign _GEN_78 = io_inputMemBlockValid ? _T_617 : inputMemBlock_77;
  assign _GEN_79 = io_inputMemBlockValid ? _T_618 : inputMemBlock_78;
  assign _GEN_80 = io_inputMemBlockValid ? _T_619 : inputMemBlock_79;
  assign _GEN_81 = io_inputMemBlockValid ? _T_620 : inputMemBlock_80;
  assign _GEN_82 = io_inputMemBlockValid ? _T_621 : inputMemBlock_81;
  assign _GEN_83 = io_inputMemBlockValid ? _T_622 : inputMemBlock_82;
  assign _GEN_84 = io_inputMemBlockValid ? _T_623 : inputMemBlock_83;
  assign _GEN_85 = io_inputMemBlockValid ? _T_624 : inputMemBlock_84;
  assign _GEN_86 = io_inputMemBlockValid ? _T_625 : inputMemBlock_85;
  assign _GEN_87 = io_inputMemBlockValid ? _T_626 : inputMemBlock_86;
  assign _GEN_88 = io_inputMemBlockValid ? _T_627 : inputMemBlock_87;
  assign _GEN_89 = io_inputMemBlockValid ? _T_628 : inputMemBlock_88;
  assign _GEN_90 = io_inputMemBlockValid ? _T_629 : inputMemBlock_89;
  assign _GEN_91 = io_inputMemBlockValid ? _T_630 : inputMemBlock_90;
  assign _GEN_92 = io_inputMemBlockValid ? _T_631 : inputMemBlock_91;
  assign _GEN_93 = io_inputMemBlockValid ? _T_632 : inputMemBlock_92;
  assign _GEN_94 = io_inputMemBlockValid ? _T_633 : inputMemBlock_93;
  assign _GEN_95 = io_inputMemBlockValid ? _T_634 : inputMemBlock_94;
  assign _GEN_96 = io_inputMemBlockValid ? _T_635 : inputMemBlock_95;
  assign _GEN_97 = io_inputMemBlockValid ? _T_636 : inputMemBlock_96;
  assign _GEN_98 = io_inputMemBlockValid ? _T_637 : inputMemBlock_97;
  assign _GEN_99 = io_inputMemBlockValid ? _T_638 : inputMemBlock_98;
  assign _GEN_100 = io_inputMemBlockValid ? _T_639 : inputMemBlock_99;
  assign _GEN_101 = io_inputMemBlockValid ? _T_640 : inputMemBlock_100;
  assign _GEN_102 = io_inputMemBlockValid ? _T_641 : inputMemBlock_101;
  assign _GEN_103 = io_inputMemBlockValid ? _T_642 : inputMemBlock_102;
  assign _GEN_104 = io_inputMemBlockValid ? _T_643 : inputMemBlock_103;
  assign _GEN_105 = io_inputMemBlockValid ? _T_644 : inputMemBlock_104;
  assign _GEN_106 = io_inputMemBlockValid ? _T_645 : inputMemBlock_105;
  assign _GEN_107 = io_inputMemBlockValid ? _T_646 : inputMemBlock_106;
  assign _GEN_108 = io_inputMemBlockValid ? _T_647 : inputMemBlock_107;
  assign _GEN_109 = io_inputMemBlockValid ? _T_648 : inputMemBlock_108;
  assign _GEN_110 = io_inputMemBlockValid ? _T_649 : inputMemBlock_109;
  assign _GEN_111 = io_inputMemBlockValid ? _T_650 : inputMemBlock_110;
  assign _GEN_112 = io_inputMemBlockValid ? _T_651 : inputMemBlock_111;
  assign _GEN_113 = io_inputMemBlockValid ? _T_652 : inputMemBlock_112;
  assign _GEN_114 = io_inputMemBlockValid ? _T_653 : inputMemBlock_113;
  assign _GEN_115 = io_inputMemBlockValid ? _T_654 : inputMemBlock_114;
  assign _GEN_116 = io_inputMemBlockValid ? _T_655 : inputMemBlock_115;
  assign _GEN_117 = io_inputMemBlockValid ? _T_656 : inputMemBlock_116;
  assign _GEN_118 = io_inputMemBlockValid ? _T_657 : inputMemBlock_117;
  assign _GEN_119 = io_inputMemBlockValid ? _T_658 : inputMemBlock_118;
  assign _GEN_120 = io_inputMemBlockValid ? _T_659 : inputMemBlock_119;
  assign _GEN_121 = io_inputMemBlockValid ? _T_660 : inputMemBlock_120;
  assign _GEN_122 = io_inputMemBlockValid ? _T_661 : inputMemBlock_121;
  assign _GEN_123 = io_inputMemBlockValid ? _T_662 : inputMemBlock_122;
  assign _GEN_124 = io_inputMemBlockValid ? _T_663 : inputMemBlock_123;
  assign _GEN_125 = io_inputMemBlockValid ? _T_664 : inputMemBlock_124;
  assign _GEN_126 = io_inputMemBlockValid ? _T_665 : inputMemBlock_125;
  assign _GEN_127 = io_inputMemBlockValid ? _T_666 : inputMemBlock_126;
  assign _GEN_128 = io_inputMemBlockValid ? _T_667 : inputMemBlock_127;
  assign _GEN_129 = io_inputMemBlockValid ? _T_668 : inputMemBlock_128;
  assign _GEN_130 = io_inputMemBlockValid ? _T_669 : inputMemBlock_129;
  assign _GEN_131 = io_inputMemBlockValid ? _T_670 : inputMemBlock_130;
  assign _GEN_132 = io_inputMemBlockValid ? _T_671 : inputMemBlock_131;
  assign _GEN_133 = io_inputMemBlockValid ? _T_672 : inputMemBlock_132;
  assign _GEN_134 = io_inputMemBlockValid ? _T_673 : inputMemBlock_133;
  assign _GEN_135 = io_inputMemBlockValid ? _T_674 : inputMemBlock_134;
  assign _GEN_136 = io_inputMemBlockValid ? _T_675 : inputMemBlock_135;
  assign _GEN_137 = io_inputMemBlockValid ? _T_676 : inputMemBlock_136;
  assign _GEN_138 = io_inputMemBlockValid ? _T_677 : inputMemBlock_137;
  assign _GEN_139 = io_inputMemBlockValid ? _T_678 : inputMemBlock_138;
  assign _GEN_140 = io_inputMemBlockValid ? _T_679 : inputMemBlock_139;
  assign _GEN_141 = io_inputMemBlockValid ? _T_680 : inputMemBlock_140;
  assign _GEN_142 = io_inputMemBlockValid ? _T_681 : inputMemBlock_141;
  assign _GEN_143 = io_inputMemBlockValid ? _T_682 : inputMemBlock_142;
  assign _GEN_144 = io_inputMemBlockValid ? _T_683 : inputMemBlock_143;
  assign _GEN_145 = io_inputMemBlockValid ? _T_684 : inputMemBlock_144;
  assign _GEN_146 = io_inputMemBlockValid ? _T_685 : inputMemBlock_145;
  assign _GEN_147 = io_inputMemBlockValid ? _T_686 : inputMemBlock_146;
  assign _GEN_148 = io_inputMemBlockValid ? _T_687 : inputMemBlock_147;
  assign _GEN_149 = io_inputMemBlockValid ? _T_688 : inputMemBlock_148;
  assign _GEN_150 = io_inputMemBlockValid ? _T_689 : inputMemBlock_149;
  assign _GEN_151 = io_inputMemBlockValid ? _T_690 : inputMemBlock_150;
  assign _GEN_152 = io_inputMemBlockValid ? _T_691 : inputMemBlock_151;
  assign _GEN_153 = io_inputMemBlockValid ? _T_692 : inputMemBlock_152;
  assign _GEN_154 = io_inputMemBlockValid ? _T_693 : inputMemBlock_153;
  assign _GEN_155 = io_inputMemBlockValid ? _T_694 : inputMemBlock_154;
  assign _GEN_156 = io_inputMemBlockValid ? _T_695 : inputMemBlock_155;
  assign _GEN_157 = io_inputMemBlockValid ? _T_696 : inputMemBlock_156;
  assign _GEN_158 = io_inputMemBlockValid ? _T_697 : inputMemBlock_157;
  assign _GEN_159 = io_inputMemBlockValid ? _T_698 : inputMemBlock_158;
  assign _GEN_160 = io_inputMemBlockValid ? _T_699 : inputMemBlock_159;
  assign _GEN_161 = io_inputMemBlockValid ? _T_700 : inputMemBlock_160;
  assign _GEN_162 = io_inputMemBlockValid ? _T_701 : inputMemBlock_161;
  assign _GEN_163 = io_inputMemBlockValid ? _T_702 : inputMemBlock_162;
  assign _GEN_164 = io_inputMemBlockValid ? _T_703 : inputMemBlock_163;
  assign _GEN_165 = io_inputMemBlockValid ? _T_704 : inputMemBlock_164;
  assign _GEN_166 = io_inputMemBlockValid ? _T_705 : inputMemBlock_165;
  assign _GEN_167 = io_inputMemBlockValid ? _T_706 : inputMemBlock_166;
  assign _GEN_168 = io_inputMemBlockValid ? _T_707 : inputMemBlock_167;
  assign _GEN_169 = io_inputMemBlockValid ? _T_708 : inputMemBlock_168;
  assign _GEN_170 = io_inputMemBlockValid ? _T_709 : inputMemBlock_169;
  assign _GEN_171 = io_inputMemBlockValid ? _T_710 : inputMemBlock_170;
  assign _GEN_172 = io_inputMemBlockValid ? _T_711 : inputMemBlock_171;
  assign _GEN_173 = io_inputMemBlockValid ? _T_712 : inputMemBlock_172;
  assign _GEN_174 = io_inputMemBlockValid ? _T_713 : inputMemBlock_173;
  assign _GEN_175 = io_inputMemBlockValid ? _T_714 : inputMemBlock_174;
  assign _GEN_176 = io_inputMemBlockValid ? _T_715 : inputMemBlock_175;
  assign _GEN_177 = io_inputMemBlockValid ? _T_716 : inputMemBlock_176;
  assign _GEN_178 = io_inputMemBlockValid ? _T_717 : inputMemBlock_177;
  assign _GEN_179 = io_inputMemBlockValid ? _T_718 : inputMemBlock_178;
  assign _GEN_180 = io_inputMemBlockValid ? _T_719 : inputMemBlock_179;
  assign _GEN_181 = io_inputMemBlockValid ? _T_720 : inputMemBlock_180;
  assign _GEN_182 = io_inputMemBlockValid ? _T_721 : inputMemBlock_181;
  assign _GEN_183 = io_inputMemBlockValid ? _T_722 : inputMemBlock_182;
  assign _GEN_184 = io_inputMemBlockValid ? _T_723 : inputMemBlock_183;
  assign _GEN_185 = io_inputMemBlockValid ? _T_724 : inputMemBlock_184;
  assign _GEN_186 = io_inputMemBlockValid ? _T_725 : inputMemBlock_185;
  assign _GEN_187 = io_inputMemBlockValid ? _T_726 : inputMemBlock_186;
  assign _GEN_188 = io_inputMemBlockValid ? _T_727 : inputMemBlock_187;
  assign _GEN_189 = io_inputMemBlockValid ? _T_728 : inputMemBlock_188;
  assign _GEN_190 = io_inputMemBlockValid ? _T_729 : inputMemBlock_189;
  assign _GEN_191 = io_inputMemBlockValid ? _T_730 : inputMemBlock_190;
  assign _GEN_192 = io_inputMemBlockValid ? _T_731 : inputMemBlock_191;
  assign _GEN_193 = io_inputMemBlockValid ? _T_732 : inputMemBlock_192;
  assign _GEN_194 = io_inputMemBlockValid ? _T_733 : inputMemBlock_193;
  assign _GEN_195 = io_inputMemBlockValid ? _T_734 : inputMemBlock_194;
  assign _GEN_196 = io_inputMemBlockValid ? _T_735 : inputMemBlock_195;
  assign _GEN_197 = io_inputMemBlockValid ? _T_736 : inputMemBlock_196;
  assign _GEN_198 = io_inputMemBlockValid ? _T_737 : inputMemBlock_197;
  assign _GEN_199 = io_inputMemBlockValid ? _T_738 : inputMemBlock_198;
  assign _GEN_200 = io_inputMemBlockValid ? _T_739 : inputMemBlock_199;
  assign _GEN_201 = io_inputMemBlockValid ? _T_740 : inputMemBlock_200;
  assign _GEN_202 = io_inputMemBlockValid ? _T_741 : inputMemBlock_201;
  assign _GEN_203 = io_inputMemBlockValid ? _T_742 : inputMemBlock_202;
  assign _GEN_204 = io_inputMemBlockValid ? _T_743 : inputMemBlock_203;
  assign _GEN_205 = io_inputMemBlockValid ? _T_744 : inputMemBlock_204;
  assign _GEN_206 = io_inputMemBlockValid ? _T_745 : inputMemBlock_205;
  assign _GEN_207 = io_inputMemBlockValid ? _T_746 : inputMemBlock_206;
  assign _GEN_208 = io_inputMemBlockValid ? _T_747 : inputMemBlock_207;
  assign _GEN_209 = io_inputMemBlockValid ? _T_748 : inputMemBlock_208;
  assign _GEN_210 = io_inputMemBlockValid ? _T_749 : inputMemBlock_209;
  assign _GEN_211 = io_inputMemBlockValid ? _T_750 : inputMemBlock_210;
  assign _GEN_212 = io_inputMemBlockValid ? _T_751 : inputMemBlock_211;
  assign _GEN_213 = io_inputMemBlockValid ? _T_752 : inputMemBlock_212;
  assign _GEN_214 = io_inputMemBlockValid ? _T_753 : inputMemBlock_213;
  assign _GEN_215 = io_inputMemBlockValid ? _T_754 : inputMemBlock_214;
  assign _GEN_216 = io_inputMemBlockValid ? _T_755 : inputMemBlock_215;
  assign _GEN_217 = io_inputMemBlockValid ? _T_756 : inputMemBlock_216;
  assign _GEN_218 = io_inputMemBlockValid ? _T_757 : inputMemBlock_217;
  assign _GEN_219 = io_inputMemBlockValid ? _T_758 : inputMemBlock_218;
  assign _GEN_220 = io_inputMemBlockValid ? _T_759 : inputMemBlock_219;
  assign _GEN_221 = io_inputMemBlockValid ? _T_760 : inputMemBlock_220;
  assign _GEN_222 = io_inputMemBlockValid ? _T_761 : inputMemBlock_221;
  assign _GEN_223 = io_inputMemBlockValid ? _T_762 : inputMemBlock_222;
  assign _GEN_224 = io_inputMemBlockValid ? _T_763 : inputMemBlock_223;
  assign _GEN_225 = io_inputMemBlockValid ? _T_764 : inputMemBlock_224;
  assign _GEN_226 = io_inputMemBlockValid ? _T_765 : inputMemBlock_225;
  assign _GEN_227 = io_inputMemBlockValid ? _T_766 : inputMemBlock_226;
  assign _GEN_228 = io_inputMemBlockValid ? _T_767 : inputMemBlock_227;
  assign _GEN_229 = io_inputMemBlockValid ? _T_768 : inputMemBlock_228;
  assign _GEN_230 = io_inputMemBlockValid ? _T_769 : inputMemBlock_229;
  assign _GEN_231 = io_inputMemBlockValid ? _T_770 : inputMemBlock_230;
  assign _GEN_232 = io_inputMemBlockValid ? _T_771 : inputMemBlock_231;
  assign _GEN_233 = io_inputMemBlockValid ? _T_772 : inputMemBlock_232;
  assign _GEN_234 = io_inputMemBlockValid ? _T_773 : inputMemBlock_233;
  assign _GEN_235 = io_inputMemBlockValid ? _T_774 : inputMemBlock_234;
  assign _GEN_236 = io_inputMemBlockValid ? _T_775 : inputMemBlock_235;
  assign _GEN_237 = io_inputMemBlockValid ? _T_776 : inputMemBlock_236;
  assign _GEN_238 = io_inputMemBlockValid ? _T_777 : inputMemBlock_237;
  assign _GEN_239 = io_inputMemBlockValid ? _T_778 : inputMemBlock_238;
  assign _GEN_240 = io_inputMemBlockValid ? _T_779 : inputMemBlock_239;
  assign _GEN_241 = io_inputMemBlockValid ? _T_780 : inputMemBlock_240;
  assign _GEN_242 = io_inputMemBlockValid ? _T_781 : inputMemBlock_241;
  assign _GEN_243 = io_inputMemBlockValid ? _T_782 : inputMemBlock_242;
  assign _GEN_244 = io_inputMemBlockValid ? _T_783 : inputMemBlock_243;
  assign _GEN_245 = io_inputMemBlockValid ? _T_784 : inputMemBlock_244;
  assign _GEN_246 = io_inputMemBlockValid ? _T_785 : inputMemBlock_245;
  assign _GEN_247 = io_inputMemBlockValid ? _T_786 : inputMemBlock_246;
  assign _GEN_248 = io_inputMemBlockValid ? _T_787 : inputMemBlock_247;
  assign _GEN_249 = io_inputMemBlockValid ? _T_788 : inputMemBlock_248;
  assign _GEN_250 = io_inputMemBlockValid ? _T_789 : inputMemBlock_249;
  assign _GEN_251 = io_inputMemBlockValid ? _T_790 : inputMemBlock_250;
  assign _GEN_252 = io_inputMemBlockValid ? _T_791 : inputMemBlock_251;
  assign _GEN_253 = io_inputMemBlockValid ? _T_792 : inputMemBlock_252;
  assign _GEN_254 = io_inputMemBlockValid ? _T_793 : inputMemBlock_253;
  assign _GEN_255 = io_inputMemBlockValid ? _T_794 : inputMemBlock_254;
  assign _GEN_256 = io_inputMemBlockValid ? _T_795 : inputMemBlock_255;
  assign _GEN_257 = io_inputMemBlockValid ? _T_796 : inputMemBlock_256;
  assign _GEN_258 = io_inputMemBlockValid ? _T_797 : inputMemBlock_257;
  assign _GEN_259 = io_inputMemBlockValid ? _T_798 : inputMemBlock_258;
  assign _GEN_260 = io_inputMemBlockValid ? _T_799 : inputMemBlock_259;
  assign _GEN_261 = io_inputMemBlockValid ? _T_800 : inputMemBlock_260;
  assign _GEN_262 = io_inputMemBlockValid ? _T_801 : inputMemBlock_261;
  assign _GEN_263 = io_inputMemBlockValid ? _T_802 : inputMemBlock_262;
  assign _GEN_264 = io_inputMemBlockValid ? _T_803 : inputMemBlock_263;
  assign _GEN_265 = io_inputMemBlockValid ? _T_804 : inputMemBlock_264;
  assign _GEN_266 = io_inputMemBlockValid ? _T_805 : inputMemBlock_265;
  assign _GEN_267 = io_inputMemBlockValid ? _T_806 : inputMemBlock_266;
  assign _GEN_268 = io_inputMemBlockValid ? _T_807 : inputMemBlock_267;
  assign _GEN_269 = io_inputMemBlockValid ? _T_808 : inputMemBlock_268;
  assign _GEN_270 = io_inputMemBlockValid ? _T_809 : inputMemBlock_269;
  assign _GEN_271 = io_inputMemBlockValid ? _T_810 : inputMemBlock_270;
  assign _GEN_272 = io_inputMemBlockValid ? _T_811 : inputMemBlock_271;
  assign _GEN_273 = io_inputMemBlockValid ? _T_812 : inputMemBlock_272;
  assign _GEN_274 = io_inputMemBlockValid ? _T_813 : inputMemBlock_273;
  assign _GEN_275 = io_inputMemBlockValid ? _T_814 : inputMemBlock_274;
  assign _GEN_276 = io_inputMemBlockValid ? _T_815 : inputMemBlock_275;
  assign _GEN_277 = io_inputMemBlockValid ? _T_816 : inputMemBlock_276;
  assign _GEN_278 = io_inputMemBlockValid ? _T_817 : inputMemBlock_277;
  assign _GEN_279 = io_inputMemBlockValid ? _T_818 : inputMemBlock_278;
  assign _GEN_280 = io_inputMemBlockValid ? _T_819 : inputMemBlock_279;
  assign _GEN_281 = io_inputMemBlockValid ? _T_820 : inputMemBlock_280;
  assign _GEN_282 = io_inputMemBlockValid ? _T_821 : inputMemBlock_281;
  assign _GEN_283 = io_inputMemBlockValid ? _T_822 : inputMemBlock_282;
  assign _GEN_284 = io_inputMemBlockValid ? _T_823 : inputMemBlock_283;
  assign _GEN_285 = io_inputMemBlockValid ? _T_824 : inputMemBlock_284;
  assign _GEN_286 = io_inputMemBlockValid ? _T_825 : inputMemBlock_285;
  assign _GEN_287 = io_inputMemBlockValid ? _T_826 : inputMemBlock_286;
  assign _GEN_288 = io_inputMemBlockValid ? _T_827 : inputMemBlock_287;
  assign _GEN_289 = io_inputMemBlockValid ? _T_828 : inputMemBlock_288;
  assign _GEN_290 = io_inputMemBlockValid ? _T_829 : inputMemBlock_289;
  assign _GEN_291 = io_inputMemBlockValid ? _T_830 : inputMemBlock_290;
  assign _GEN_292 = io_inputMemBlockValid ? _T_831 : inputMemBlock_291;
  assign _GEN_293 = io_inputMemBlockValid ? _T_832 : inputMemBlock_292;
  assign _GEN_294 = io_inputMemBlockValid ? _T_833 : inputMemBlock_293;
  assign _GEN_295 = io_inputMemBlockValid ? _T_834 : inputMemBlock_294;
  assign _GEN_296 = io_inputMemBlockValid ? _T_835 : inputMemBlock_295;
  assign _GEN_297 = io_inputMemBlockValid ? _T_836 : inputMemBlock_296;
  assign _GEN_298 = io_inputMemBlockValid ? _T_837 : inputMemBlock_297;
  assign _GEN_299 = io_inputMemBlockValid ? _T_838 : inputMemBlock_298;
  assign _GEN_300 = io_inputMemBlockValid ? _T_839 : inputMemBlock_299;
  assign _GEN_301 = io_inputMemBlockValid ? _T_840 : inputMemBlock_300;
  assign _GEN_302 = io_inputMemBlockValid ? _T_841 : inputMemBlock_301;
  assign _GEN_303 = io_inputMemBlockValid ? _T_842 : inputMemBlock_302;
  assign _GEN_304 = io_inputMemBlockValid ? _T_843 : inputMemBlock_303;
  assign _GEN_305 = io_inputMemBlockValid ? _T_844 : inputMemBlock_304;
  assign _GEN_306 = io_inputMemBlockValid ? _T_845 : inputMemBlock_305;
  assign _GEN_307 = io_inputMemBlockValid ? _T_846 : inputMemBlock_306;
  assign _GEN_308 = io_inputMemBlockValid ? _T_847 : inputMemBlock_307;
  assign _GEN_309 = io_inputMemBlockValid ? _T_848 : inputMemBlock_308;
  assign _GEN_310 = io_inputMemBlockValid ? _T_849 : inputMemBlock_309;
  assign _GEN_311 = io_inputMemBlockValid ? _T_850 : inputMemBlock_310;
  assign _GEN_312 = io_inputMemBlockValid ? _T_851 : inputMemBlock_311;
  assign _GEN_313 = io_inputMemBlockValid ? _T_852 : inputMemBlock_312;
  assign _GEN_314 = io_inputMemBlockValid ? _T_853 : inputMemBlock_313;
  assign _GEN_315 = io_inputMemBlockValid ? _T_854 : inputMemBlock_314;
  assign _GEN_316 = io_inputMemBlockValid ? _T_855 : inputMemBlock_315;
  assign _GEN_317 = io_inputMemBlockValid ? _T_856 : inputMemBlock_316;
  assign _GEN_318 = io_inputMemBlockValid ? _T_857 : inputMemBlock_317;
  assign _GEN_319 = io_inputMemBlockValid ? _T_858 : inputMemBlock_318;
  assign _GEN_320 = io_inputMemBlockValid ? _T_859 : inputMemBlock_319;
  assign _GEN_321 = io_inputMemBlockValid ? _T_860 : inputMemBlock_320;
  assign _GEN_322 = io_inputMemBlockValid ? _T_861 : inputMemBlock_321;
  assign _GEN_323 = io_inputMemBlockValid ? _T_862 : inputMemBlock_322;
  assign _GEN_324 = io_inputMemBlockValid ? _T_863 : inputMemBlock_323;
  assign _GEN_325 = io_inputMemBlockValid ? _T_864 : inputMemBlock_324;
  assign _GEN_326 = io_inputMemBlockValid ? _T_865 : inputMemBlock_325;
  assign _GEN_327 = io_inputMemBlockValid ? _T_866 : inputMemBlock_326;
  assign _GEN_328 = io_inputMemBlockValid ? _T_867 : inputMemBlock_327;
  assign _GEN_329 = io_inputMemBlockValid ? _T_868 : inputMemBlock_328;
  assign _GEN_330 = io_inputMemBlockValid ? _T_869 : inputMemBlock_329;
  assign _GEN_331 = io_inputMemBlockValid ? _T_870 : inputMemBlock_330;
  assign _GEN_332 = io_inputMemBlockValid ? _T_871 : inputMemBlock_331;
  assign _GEN_333 = io_inputMemBlockValid ? _T_872 : inputMemBlock_332;
  assign _GEN_334 = io_inputMemBlockValid ? _T_873 : inputMemBlock_333;
  assign _GEN_335 = io_inputMemBlockValid ? _T_874 : inputMemBlock_334;
  assign _GEN_336 = io_inputMemBlockValid ? _T_875 : inputMemBlock_335;
  assign _GEN_337 = io_inputMemBlockValid ? _T_876 : inputMemBlock_336;
  assign _GEN_338 = io_inputMemBlockValid ? _T_877 : inputMemBlock_337;
  assign _GEN_339 = io_inputMemBlockValid ? _T_878 : inputMemBlock_338;
  assign _GEN_340 = io_inputMemBlockValid ? _T_879 : inputMemBlock_339;
  assign _GEN_341 = io_inputMemBlockValid ? _T_880 : inputMemBlock_340;
  assign _GEN_342 = io_inputMemBlockValid ? _T_881 : inputMemBlock_341;
  assign _GEN_343 = io_inputMemBlockValid ? _T_882 : inputMemBlock_342;
  assign _GEN_344 = io_inputMemBlockValid ? _T_883 : inputMemBlock_343;
  assign _GEN_345 = io_inputMemBlockValid ? _T_884 : inputMemBlock_344;
  assign _GEN_346 = io_inputMemBlockValid ? _T_885 : inputMemBlock_345;
  assign _GEN_347 = io_inputMemBlockValid ? _T_886 : inputMemBlock_346;
  assign _GEN_348 = io_inputMemBlockValid ? _T_887 : inputMemBlock_347;
  assign _GEN_349 = io_inputMemBlockValid ? _T_888 : inputMemBlock_348;
  assign _GEN_350 = io_inputMemBlockValid ? _T_889 : inputMemBlock_349;
  assign _GEN_351 = io_inputMemBlockValid ? _T_890 : inputMemBlock_350;
  assign _GEN_352 = io_inputMemBlockValid ? _T_891 : inputMemBlock_351;
  assign _GEN_353 = io_inputMemBlockValid ? _T_892 : inputMemBlock_352;
  assign _GEN_354 = io_inputMemBlockValid ? _T_893 : inputMemBlock_353;
  assign _GEN_355 = io_inputMemBlockValid ? _T_894 : inputMemBlock_354;
  assign _GEN_356 = io_inputMemBlockValid ? _T_895 : inputMemBlock_355;
  assign _GEN_357 = io_inputMemBlockValid ? _T_896 : inputMemBlock_356;
  assign _GEN_358 = io_inputMemBlockValid ? _T_897 : inputMemBlock_357;
  assign _GEN_359 = io_inputMemBlockValid ? _T_898 : inputMemBlock_358;
  assign _GEN_360 = io_inputMemBlockValid ? _T_899 : inputMemBlock_359;
  assign _GEN_361 = io_inputMemBlockValid ? _T_900 : inputMemBlock_360;
  assign _GEN_362 = io_inputMemBlockValid ? _T_901 : inputMemBlock_361;
  assign _GEN_363 = io_inputMemBlockValid ? _T_902 : inputMemBlock_362;
  assign _GEN_364 = io_inputMemBlockValid ? _T_903 : inputMemBlock_363;
  assign _GEN_365 = io_inputMemBlockValid ? _T_904 : inputMemBlock_364;
  assign _GEN_366 = io_inputMemBlockValid ? _T_905 : inputMemBlock_365;
  assign _GEN_367 = io_inputMemBlockValid ? _T_906 : inputMemBlock_366;
  assign _GEN_368 = io_inputMemBlockValid ? _T_907 : inputMemBlock_367;
  assign _GEN_369 = io_inputMemBlockValid ? _T_908 : inputMemBlock_368;
  assign _GEN_370 = io_inputMemBlockValid ? _T_909 : inputMemBlock_369;
  assign _GEN_371 = io_inputMemBlockValid ? _T_910 : inputMemBlock_370;
  assign _GEN_372 = io_inputMemBlockValid ? _T_911 : inputMemBlock_371;
  assign _GEN_373 = io_inputMemBlockValid ? _T_912 : inputMemBlock_372;
  assign _GEN_374 = io_inputMemBlockValid ? _T_913 : inputMemBlock_373;
  assign _GEN_375 = io_inputMemBlockValid ? _T_914 : inputMemBlock_374;
  assign _GEN_376 = io_inputMemBlockValid ? _T_915 : inputMemBlock_375;
  assign _GEN_377 = io_inputMemBlockValid ? _T_916 : inputMemBlock_376;
  assign _GEN_378 = io_inputMemBlockValid ? _T_917 : inputMemBlock_377;
  assign _GEN_379 = io_inputMemBlockValid ? _T_918 : inputMemBlock_378;
  assign _GEN_380 = io_inputMemBlockValid ? _T_919 : inputMemBlock_379;
  assign _GEN_381 = io_inputMemBlockValid ? _T_920 : inputMemBlock_380;
  assign _GEN_382 = io_inputMemBlockValid ? _T_921 : inputMemBlock_381;
  assign _GEN_383 = io_inputMemBlockValid ? _T_922 : inputMemBlock_382;
  assign _GEN_384 = io_inputMemBlockValid ? _T_923 : inputMemBlock_383;
  assign _GEN_385 = io_inputMemBlockValid ? _T_924 : inputMemBlock_384;
  assign _GEN_386 = io_inputMemBlockValid ? _T_925 : inputMemBlock_385;
  assign _GEN_387 = io_inputMemBlockValid ? _T_926 : inputMemBlock_386;
  assign _GEN_388 = io_inputMemBlockValid ? _T_927 : inputMemBlock_387;
  assign _GEN_389 = io_inputMemBlockValid ? _T_928 : inputMemBlock_388;
  assign _GEN_390 = io_inputMemBlockValid ? _T_929 : inputMemBlock_389;
  assign _GEN_391 = io_inputMemBlockValid ? _T_930 : inputMemBlock_390;
  assign _GEN_392 = io_inputMemBlockValid ? _T_931 : inputMemBlock_391;
  assign _GEN_393 = io_inputMemBlockValid ? _T_932 : inputMemBlock_392;
  assign _GEN_394 = io_inputMemBlockValid ? _T_933 : inputMemBlock_393;
  assign _GEN_395 = io_inputMemBlockValid ? _T_934 : inputMemBlock_394;
  assign _GEN_396 = io_inputMemBlockValid ? _T_935 : inputMemBlock_395;
  assign _GEN_397 = io_inputMemBlockValid ? _T_936 : inputMemBlock_396;
  assign _GEN_398 = io_inputMemBlockValid ? _T_937 : inputMemBlock_397;
  assign _GEN_399 = io_inputMemBlockValid ? _T_938 : inputMemBlock_398;
  assign _GEN_400 = io_inputMemBlockValid ? _T_939 : inputMemBlock_399;
  assign _GEN_401 = io_inputMemBlockValid ? _T_940 : inputMemBlock_400;
  assign _GEN_402 = io_inputMemBlockValid ? _T_941 : inputMemBlock_401;
  assign _GEN_403 = io_inputMemBlockValid ? _T_942 : inputMemBlock_402;
  assign _GEN_404 = io_inputMemBlockValid ? _T_943 : inputMemBlock_403;
  assign _GEN_405 = io_inputMemBlockValid ? _T_944 : inputMemBlock_404;
  assign _GEN_406 = io_inputMemBlockValid ? _T_945 : inputMemBlock_405;
  assign _GEN_407 = io_inputMemBlockValid ? _T_946 : inputMemBlock_406;
  assign _GEN_408 = io_inputMemBlockValid ? _T_947 : inputMemBlock_407;
  assign _GEN_409 = io_inputMemBlockValid ? _T_948 : inputMemBlock_408;
  assign _GEN_410 = io_inputMemBlockValid ? _T_949 : inputMemBlock_409;
  assign _GEN_411 = io_inputMemBlockValid ? _T_950 : inputMemBlock_410;
  assign _GEN_412 = io_inputMemBlockValid ? _T_951 : inputMemBlock_411;
  assign _GEN_413 = io_inputMemBlockValid ? _T_952 : inputMemBlock_412;
  assign _GEN_414 = io_inputMemBlockValid ? _T_953 : inputMemBlock_413;
  assign _GEN_415 = io_inputMemBlockValid ? _T_954 : inputMemBlock_414;
  assign _GEN_416 = io_inputMemBlockValid ? _T_955 : inputMemBlock_415;
  assign _GEN_417 = io_inputMemBlockValid ? _T_956 : inputMemBlock_416;
  assign _GEN_418 = io_inputMemBlockValid ? _T_957 : inputMemBlock_417;
  assign _GEN_419 = io_inputMemBlockValid ? _T_958 : inputMemBlock_418;
  assign _GEN_420 = io_inputMemBlockValid ? _T_959 : inputMemBlock_419;
  assign _GEN_421 = io_inputMemBlockValid ? _T_960 : inputMemBlock_420;
  assign _GEN_422 = io_inputMemBlockValid ? _T_961 : inputMemBlock_421;
  assign _GEN_423 = io_inputMemBlockValid ? _T_962 : inputMemBlock_422;
  assign _GEN_424 = io_inputMemBlockValid ? _T_963 : inputMemBlock_423;
  assign _GEN_425 = io_inputMemBlockValid ? _T_964 : inputMemBlock_424;
  assign _GEN_426 = io_inputMemBlockValid ? _T_965 : inputMemBlock_425;
  assign _GEN_427 = io_inputMemBlockValid ? _T_966 : inputMemBlock_426;
  assign _GEN_428 = io_inputMemBlockValid ? _T_967 : inputMemBlock_427;
  assign _GEN_429 = io_inputMemBlockValid ? _T_968 : inputMemBlock_428;
  assign _GEN_430 = io_inputMemBlockValid ? _T_969 : inputMemBlock_429;
  assign _GEN_431 = io_inputMemBlockValid ? _T_970 : inputMemBlock_430;
  assign _GEN_432 = io_inputMemBlockValid ? _T_971 : inputMemBlock_431;
  assign _GEN_433 = io_inputMemBlockValid ? _T_972 : inputMemBlock_432;
  assign _GEN_434 = io_inputMemBlockValid ? _T_973 : inputMemBlock_433;
  assign _GEN_435 = io_inputMemBlockValid ? _T_974 : inputMemBlock_434;
  assign _GEN_436 = io_inputMemBlockValid ? _T_975 : inputMemBlock_435;
  assign _GEN_437 = io_inputMemBlockValid ? _T_976 : inputMemBlock_436;
  assign _GEN_438 = io_inputMemBlockValid ? _T_977 : inputMemBlock_437;
  assign _GEN_439 = io_inputMemBlockValid ? _T_978 : inputMemBlock_438;
  assign _GEN_440 = io_inputMemBlockValid ? _T_979 : inputMemBlock_439;
  assign _GEN_441 = io_inputMemBlockValid ? _T_980 : inputMemBlock_440;
  assign _GEN_442 = io_inputMemBlockValid ? _T_981 : inputMemBlock_441;
  assign _GEN_443 = io_inputMemBlockValid ? _T_982 : inputMemBlock_442;
  assign _GEN_444 = io_inputMemBlockValid ? _T_983 : inputMemBlock_443;
  assign _GEN_445 = io_inputMemBlockValid ? _T_984 : inputMemBlock_444;
  assign _GEN_446 = io_inputMemBlockValid ? _T_985 : inputMemBlock_445;
  assign _GEN_447 = io_inputMemBlockValid ? _T_986 : inputMemBlock_446;
  assign _GEN_448 = io_inputMemBlockValid ? _T_987 : inputMemBlock_447;
  assign _GEN_449 = io_inputMemBlockValid ? _T_988 : inputMemBlock_448;
  assign _GEN_450 = io_inputMemBlockValid ? _T_989 : inputMemBlock_449;
  assign _GEN_451 = io_inputMemBlockValid ? _T_990 : inputMemBlock_450;
  assign _GEN_452 = io_inputMemBlockValid ? _T_991 : inputMemBlock_451;
  assign _GEN_453 = io_inputMemBlockValid ? _T_992 : inputMemBlock_452;
  assign _GEN_454 = io_inputMemBlockValid ? _T_993 : inputMemBlock_453;
  assign _GEN_455 = io_inputMemBlockValid ? _T_994 : inputMemBlock_454;
  assign _GEN_456 = io_inputMemBlockValid ? _T_995 : inputMemBlock_455;
  assign _GEN_457 = io_inputMemBlockValid ? _T_996 : inputMemBlock_456;
  assign _GEN_458 = io_inputMemBlockValid ? _T_997 : inputMemBlock_457;
  assign _GEN_459 = io_inputMemBlockValid ? _T_998 : inputMemBlock_458;
  assign _GEN_460 = io_inputMemBlockValid ? _T_999 : inputMemBlock_459;
  assign _GEN_461 = io_inputMemBlockValid ? _T_1000 : inputMemBlock_460;
  assign _GEN_462 = io_inputMemBlockValid ? _T_1001 : inputMemBlock_461;
  assign _GEN_463 = io_inputMemBlockValid ? _T_1002 : inputMemBlock_462;
  assign _GEN_464 = io_inputMemBlockValid ? _T_1003 : inputMemBlock_463;
  assign _GEN_465 = io_inputMemBlockValid ? _T_1004 : inputMemBlock_464;
  assign _GEN_466 = io_inputMemBlockValid ? _T_1005 : inputMemBlock_465;
  assign _GEN_467 = io_inputMemBlockValid ? _T_1006 : inputMemBlock_466;
  assign _GEN_468 = io_inputMemBlockValid ? _T_1007 : inputMemBlock_467;
  assign _GEN_469 = io_inputMemBlockValid ? _T_1008 : inputMemBlock_468;
  assign _GEN_470 = io_inputMemBlockValid ? _T_1009 : inputMemBlock_469;
  assign _GEN_471 = io_inputMemBlockValid ? _T_1010 : inputMemBlock_470;
  assign _GEN_472 = io_inputMemBlockValid ? _T_1011 : inputMemBlock_471;
  assign _GEN_473 = io_inputMemBlockValid ? _T_1012 : inputMemBlock_472;
  assign _GEN_474 = io_inputMemBlockValid ? _T_1013 : inputMemBlock_473;
  assign _GEN_475 = io_inputMemBlockValid ? _T_1014 : inputMemBlock_474;
  assign _GEN_476 = io_inputMemBlockValid ? _T_1015 : inputMemBlock_475;
  assign _GEN_477 = io_inputMemBlockValid ? _T_1016 : inputMemBlock_476;
  assign _GEN_478 = io_inputMemBlockValid ? _T_1017 : inputMemBlock_477;
  assign _GEN_479 = io_inputMemBlockValid ? _T_1018 : inputMemBlock_478;
  assign _GEN_480 = io_inputMemBlockValid ? _T_1019 : inputMemBlock_479;
  assign _GEN_481 = io_inputMemBlockValid ? _T_1020 : inputMemBlock_480;
  assign _GEN_482 = io_inputMemBlockValid ? _T_1021 : inputMemBlock_481;
  assign _GEN_483 = io_inputMemBlockValid ? _T_1022 : inputMemBlock_482;
  assign _GEN_484 = io_inputMemBlockValid ? _T_1023 : inputMemBlock_483;
  assign _GEN_485 = io_inputMemBlockValid ? _T_1024 : inputMemBlock_484;
  assign _GEN_486 = io_inputMemBlockValid ? _T_1025 : inputMemBlock_485;
  assign _GEN_487 = io_inputMemBlockValid ? _T_1026 : inputMemBlock_486;
  assign _GEN_488 = io_inputMemBlockValid ? _T_1027 : inputMemBlock_487;
  assign _GEN_489 = io_inputMemBlockValid ? _T_1028 : inputMemBlock_488;
  assign _GEN_490 = io_inputMemBlockValid ? _T_1029 : inputMemBlock_489;
  assign _GEN_491 = io_inputMemBlockValid ? _T_1030 : inputMemBlock_490;
  assign _GEN_492 = io_inputMemBlockValid ? _T_1031 : inputMemBlock_491;
  assign _GEN_493 = io_inputMemBlockValid ? _T_1032 : inputMemBlock_492;
  assign _GEN_494 = io_inputMemBlockValid ? _T_1033 : inputMemBlock_493;
  assign _GEN_495 = io_inputMemBlockValid ? _T_1034 : inputMemBlock_494;
  assign _GEN_496 = io_inputMemBlockValid ? _T_1035 : inputMemBlock_495;
  assign _GEN_497 = io_inputMemBlockValid ? _T_1036 : inputMemBlock_496;
  assign _GEN_498 = io_inputMemBlockValid ? _T_1037 : inputMemBlock_497;
  assign _GEN_499 = io_inputMemBlockValid ? _T_1038 : inputMemBlock_498;
  assign _GEN_500 = io_inputMemBlockValid ? _T_1039 : inputMemBlock_499;
  assign _GEN_501 = io_inputMemBlockValid ? _T_1040 : inputMemBlock_500;
  assign _GEN_502 = io_inputMemBlockValid ? _T_1041 : inputMemBlock_501;
  assign _GEN_503 = io_inputMemBlockValid ? _T_1042 : inputMemBlock_502;
  assign _GEN_504 = io_inputMemBlockValid ? _T_1043 : inputMemBlock_503;
  assign _GEN_505 = io_inputMemBlockValid ? _T_1044 : inputMemBlock_504;
  assign _GEN_506 = io_inputMemBlockValid ? _T_1045 : inputMemBlock_505;
  assign _GEN_507 = io_inputMemBlockValid ? _T_1046 : inputMemBlock_506;
  assign _GEN_508 = io_inputMemBlockValid ? _T_1047 : inputMemBlock_507;
  assign _GEN_509 = io_inputMemBlockValid ? _T_1048 : inputMemBlock_508;
  assign _GEN_510 = io_inputMemBlockValid ? _T_1049 : inputMemBlock_509;
  assign _GEN_511 = io_inputMemBlockValid ? _T_1050 : inputMemBlock_510;
  assign _GEN_512 = io_inputMemBlockValid ? _T_1051 : inputMemBlock_511;
  assign _T_1053 = inputBitsRemaining == 10'h0;
  assign _T_1055 = io_inputFinished == 1'h0;
  assign _T_1056 = _T_1053 & _T_1055;
  assign nextBitValid = inputAdvance;
  assign nextBit = inputMemBlock_0;
  assign inputAdvance = _T_1582;
  assign _T_1579 = outputBits != 10'h200;
  assign _T_1581 = inputBitsRemaining != 10'h0;
  assign _T_1582 = _T_1579 & _T_1581;
  assign _T_1584 = inputBitsRemaining - 10'h1;
  assign _T_1585 = _T_1584[9:0];
  assign _GEN_513 = inputAdvance ? _T_1585 : _GEN_0;
  assign _GEN_514 = inputAdvance ? inputMemBlock_1 : _GEN_1;
  assign _GEN_515 = inputAdvance ? inputMemBlock_2 : _GEN_2;
  assign _GEN_516 = inputAdvance ? inputMemBlock_3 : _GEN_3;
  assign _GEN_517 = inputAdvance ? inputMemBlock_4 : _GEN_4;
  assign _GEN_518 = inputAdvance ? inputMemBlock_5 : _GEN_5;
  assign _GEN_519 = inputAdvance ? inputMemBlock_6 : _GEN_6;
  assign _GEN_520 = inputAdvance ? inputMemBlock_7 : _GEN_7;
  assign _GEN_521 = inputAdvance ? inputMemBlock_8 : _GEN_8;
  assign _GEN_522 = inputAdvance ? inputMemBlock_9 : _GEN_9;
  assign _GEN_523 = inputAdvance ? inputMemBlock_10 : _GEN_10;
  assign _GEN_524 = inputAdvance ? inputMemBlock_11 : _GEN_11;
  assign _GEN_525 = inputAdvance ? inputMemBlock_12 : _GEN_12;
  assign _GEN_526 = inputAdvance ? inputMemBlock_13 : _GEN_13;
  assign _GEN_527 = inputAdvance ? inputMemBlock_14 : _GEN_14;
  assign _GEN_528 = inputAdvance ? inputMemBlock_15 : _GEN_15;
  assign _GEN_529 = inputAdvance ? inputMemBlock_16 : _GEN_16;
  assign _GEN_530 = inputAdvance ? inputMemBlock_17 : _GEN_17;
  assign _GEN_531 = inputAdvance ? inputMemBlock_18 : _GEN_18;
  assign _GEN_532 = inputAdvance ? inputMemBlock_19 : _GEN_19;
  assign _GEN_533 = inputAdvance ? inputMemBlock_20 : _GEN_20;
  assign _GEN_534 = inputAdvance ? inputMemBlock_21 : _GEN_21;
  assign _GEN_535 = inputAdvance ? inputMemBlock_22 : _GEN_22;
  assign _GEN_536 = inputAdvance ? inputMemBlock_23 : _GEN_23;
  assign _GEN_537 = inputAdvance ? inputMemBlock_24 : _GEN_24;
  assign _GEN_538 = inputAdvance ? inputMemBlock_25 : _GEN_25;
  assign _GEN_539 = inputAdvance ? inputMemBlock_26 : _GEN_26;
  assign _GEN_540 = inputAdvance ? inputMemBlock_27 : _GEN_27;
  assign _GEN_541 = inputAdvance ? inputMemBlock_28 : _GEN_28;
  assign _GEN_542 = inputAdvance ? inputMemBlock_29 : _GEN_29;
  assign _GEN_543 = inputAdvance ? inputMemBlock_30 : _GEN_30;
  assign _GEN_544 = inputAdvance ? inputMemBlock_31 : _GEN_31;
  assign _GEN_545 = inputAdvance ? inputMemBlock_32 : _GEN_32;
  assign _GEN_546 = inputAdvance ? inputMemBlock_33 : _GEN_33;
  assign _GEN_547 = inputAdvance ? inputMemBlock_34 : _GEN_34;
  assign _GEN_548 = inputAdvance ? inputMemBlock_35 : _GEN_35;
  assign _GEN_549 = inputAdvance ? inputMemBlock_36 : _GEN_36;
  assign _GEN_550 = inputAdvance ? inputMemBlock_37 : _GEN_37;
  assign _GEN_551 = inputAdvance ? inputMemBlock_38 : _GEN_38;
  assign _GEN_552 = inputAdvance ? inputMemBlock_39 : _GEN_39;
  assign _GEN_553 = inputAdvance ? inputMemBlock_40 : _GEN_40;
  assign _GEN_554 = inputAdvance ? inputMemBlock_41 : _GEN_41;
  assign _GEN_555 = inputAdvance ? inputMemBlock_42 : _GEN_42;
  assign _GEN_556 = inputAdvance ? inputMemBlock_43 : _GEN_43;
  assign _GEN_557 = inputAdvance ? inputMemBlock_44 : _GEN_44;
  assign _GEN_558 = inputAdvance ? inputMemBlock_45 : _GEN_45;
  assign _GEN_559 = inputAdvance ? inputMemBlock_46 : _GEN_46;
  assign _GEN_560 = inputAdvance ? inputMemBlock_47 : _GEN_47;
  assign _GEN_561 = inputAdvance ? inputMemBlock_48 : _GEN_48;
  assign _GEN_562 = inputAdvance ? inputMemBlock_49 : _GEN_49;
  assign _GEN_563 = inputAdvance ? inputMemBlock_50 : _GEN_50;
  assign _GEN_564 = inputAdvance ? inputMemBlock_51 : _GEN_51;
  assign _GEN_565 = inputAdvance ? inputMemBlock_52 : _GEN_52;
  assign _GEN_566 = inputAdvance ? inputMemBlock_53 : _GEN_53;
  assign _GEN_567 = inputAdvance ? inputMemBlock_54 : _GEN_54;
  assign _GEN_568 = inputAdvance ? inputMemBlock_55 : _GEN_55;
  assign _GEN_569 = inputAdvance ? inputMemBlock_56 : _GEN_56;
  assign _GEN_570 = inputAdvance ? inputMemBlock_57 : _GEN_57;
  assign _GEN_571 = inputAdvance ? inputMemBlock_58 : _GEN_58;
  assign _GEN_572 = inputAdvance ? inputMemBlock_59 : _GEN_59;
  assign _GEN_573 = inputAdvance ? inputMemBlock_60 : _GEN_60;
  assign _GEN_574 = inputAdvance ? inputMemBlock_61 : _GEN_61;
  assign _GEN_575 = inputAdvance ? inputMemBlock_62 : _GEN_62;
  assign _GEN_576 = inputAdvance ? inputMemBlock_63 : _GEN_63;
  assign _GEN_577 = inputAdvance ? inputMemBlock_64 : _GEN_64;
  assign _GEN_578 = inputAdvance ? inputMemBlock_65 : _GEN_65;
  assign _GEN_579 = inputAdvance ? inputMemBlock_66 : _GEN_66;
  assign _GEN_580 = inputAdvance ? inputMemBlock_67 : _GEN_67;
  assign _GEN_581 = inputAdvance ? inputMemBlock_68 : _GEN_68;
  assign _GEN_582 = inputAdvance ? inputMemBlock_69 : _GEN_69;
  assign _GEN_583 = inputAdvance ? inputMemBlock_70 : _GEN_70;
  assign _GEN_584 = inputAdvance ? inputMemBlock_71 : _GEN_71;
  assign _GEN_585 = inputAdvance ? inputMemBlock_72 : _GEN_72;
  assign _GEN_586 = inputAdvance ? inputMemBlock_73 : _GEN_73;
  assign _GEN_587 = inputAdvance ? inputMemBlock_74 : _GEN_74;
  assign _GEN_588 = inputAdvance ? inputMemBlock_75 : _GEN_75;
  assign _GEN_589 = inputAdvance ? inputMemBlock_76 : _GEN_76;
  assign _GEN_590 = inputAdvance ? inputMemBlock_77 : _GEN_77;
  assign _GEN_591 = inputAdvance ? inputMemBlock_78 : _GEN_78;
  assign _GEN_592 = inputAdvance ? inputMemBlock_79 : _GEN_79;
  assign _GEN_593 = inputAdvance ? inputMemBlock_80 : _GEN_80;
  assign _GEN_594 = inputAdvance ? inputMemBlock_81 : _GEN_81;
  assign _GEN_595 = inputAdvance ? inputMemBlock_82 : _GEN_82;
  assign _GEN_596 = inputAdvance ? inputMemBlock_83 : _GEN_83;
  assign _GEN_597 = inputAdvance ? inputMemBlock_84 : _GEN_84;
  assign _GEN_598 = inputAdvance ? inputMemBlock_85 : _GEN_85;
  assign _GEN_599 = inputAdvance ? inputMemBlock_86 : _GEN_86;
  assign _GEN_600 = inputAdvance ? inputMemBlock_87 : _GEN_87;
  assign _GEN_601 = inputAdvance ? inputMemBlock_88 : _GEN_88;
  assign _GEN_602 = inputAdvance ? inputMemBlock_89 : _GEN_89;
  assign _GEN_603 = inputAdvance ? inputMemBlock_90 : _GEN_90;
  assign _GEN_604 = inputAdvance ? inputMemBlock_91 : _GEN_91;
  assign _GEN_605 = inputAdvance ? inputMemBlock_92 : _GEN_92;
  assign _GEN_606 = inputAdvance ? inputMemBlock_93 : _GEN_93;
  assign _GEN_607 = inputAdvance ? inputMemBlock_94 : _GEN_94;
  assign _GEN_608 = inputAdvance ? inputMemBlock_95 : _GEN_95;
  assign _GEN_609 = inputAdvance ? inputMemBlock_96 : _GEN_96;
  assign _GEN_610 = inputAdvance ? inputMemBlock_97 : _GEN_97;
  assign _GEN_611 = inputAdvance ? inputMemBlock_98 : _GEN_98;
  assign _GEN_612 = inputAdvance ? inputMemBlock_99 : _GEN_99;
  assign _GEN_613 = inputAdvance ? inputMemBlock_100 : _GEN_100;
  assign _GEN_614 = inputAdvance ? inputMemBlock_101 : _GEN_101;
  assign _GEN_615 = inputAdvance ? inputMemBlock_102 : _GEN_102;
  assign _GEN_616 = inputAdvance ? inputMemBlock_103 : _GEN_103;
  assign _GEN_617 = inputAdvance ? inputMemBlock_104 : _GEN_104;
  assign _GEN_618 = inputAdvance ? inputMemBlock_105 : _GEN_105;
  assign _GEN_619 = inputAdvance ? inputMemBlock_106 : _GEN_106;
  assign _GEN_620 = inputAdvance ? inputMemBlock_107 : _GEN_107;
  assign _GEN_621 = inputAdvance ? inputMemBlock_108 : _GEN_108;
  assign _GEN_622 = inputAdvance ? inputMemBlock_109 : _GEN_109;
  assign _GEN_623 = inputAdvance ? inputMemBlock_110 : _GEN_110;
  assign _GEN_624 = inputAdvance ? inputMemBlock_111 : _GEN_111;
  assign _GEN_625 = inputAdvance ? inputMemBlock_112 : _GEN_112;
  assign _GEN_626 = inputAdvance ? inputMemBlock_113 : _GEN_113;
  assign _GEN_627 = inputAdvance ? inputMemBlock_114 : _GEN_114;
  assign _GEN_628 = inputAdvance ? inputMemBlock_115 : _GEN_115;
  assign _GEN_629 = inputAdvance ? inputMemBlock_116 : _GEN_116;
  assign _GEN_630 = inputAdvance ? inputMemBlock_117 : _GEN_117;
  assign _GEN_631 = inputAdvance ? inputMemBlock_118 : _GEN_118;
  assign _GEN_632 = inputAdvance ? inputMemBlock_119 : _GEN_119;
  assign _GEN_633 = inputAdvance ? inputMemBlock_120 : _GEN_120;
  assign _GEN_634 = inputAdvance ? inputMemBlock_121 : _GEN_121;
  assign _GEN_635 = inputAdvance ? inputMemBlock_122 : _GEN_122;
  assign _GEN_636 = inputAdvance ? inputMemBlock_123 : _GEN_123;
  assign _GEN_637 = inputAdvance ? inputMemBlock_124 : _GEN_124;
  assign _GEN_638 = inputAdvance ? inputMemBlock_125 : _GEN_125;
  assign _GEN_639 = inputAdvance ? inputMemBlock_126 : _GEN_126;
  assign _GEN_640 = inputAdvance ? inputMemBlock_127 : _GEN_127;
  assign _GEN_641 = inputAdvance ? inputMemBlock_128 : _GEN_128;
  assign _GEN_642 = inputAdvance ? inputMemBlock_129 : _GEN_129;
  assign _GEN_643 = inputAdvance ? inputMemBlock_130 : _GEN_130;
  assign _GEN_644 = inputAdvance ? inputMemBlock_131 : _GEN_131;
  assign _GEN_645 = inputAdvance ? inputMemBlock_132 : _GEN_132;
  assign _GEN_646 = inputAdvance ? inputMemBlock_133 : _GEN_133;
  assign _GEN_647 = inputAdvance ? inputMemBlock_134 : _GEN_134;
  assign _GEN_648 = inputAdvance ? inputMemBlock_135 : _GEN_135;
  assign _GEN_649 = inputAdvance ? inputMemBlock_136 : _GEN_136;
  assign _GEN_650 = inputAdvance ? inputMemBlock_137 : _GEN_137;
  assign _GEN_651 = inputAdvance ? inputMemBlock_138 : _GEN_138;
  assign _GEN_652 = inputAdvance ? inputMemBlock_139 : _GEN_139;
  assign _GEN_653 = inputAdvance ? inputMemBlock_140 : _GEN_140;
  assign _GEN_654 = inputAdvance ? inputMemBlock_141 : _GEN_141;
  assign _GEN_655 = inputAdvance ? inputMemBlock_142 : _GEN_142;
  assign _GEN_656 = inputAdvance ? inputMemBlock_143 : _GEN_143;
  assign _GEN_657 = inputAdvance ? inputMemBlock_144 : _GEN_144;
  assign _GEN_658 = inputAdvance ? inputMemBlock_145 : _GEN_145;
  assign _GEN_659 = inputAdvance ? inputMemBlock_146 : _GEN_146;
  assign _GEN_660 = inputAdvance ? inputMemBlock_147 : _GEN_147;
  assign _GEN_661 = inputAdvance ? inputMemBlock_148 : _GEN_148;
  assign _GEN_662 = inputAdvance ? inputMemBlock_149 : _GEN_149;
  assign _GEN_663 = inputAdvance ? inputMemBlock_150 : _GEN_150;
  assign _GEN_664 = inputAdvance ? inputMemBlock_151 : _GEN_151;
  assign _GEN_665 = inputAdvance ? inputMemBlock_152 : _GEN_152;
  assign _GEN_666 = inputAdvance ? inputMemBlock_153 : _GEN_153;
  assign _GEN_667 = inputAdvance ? inputMemBlock_154 : _GEN_154;
  assign _GEN_668 = inputAdvance ? inputMemBlock_155 : _GEN_155;
  assign _GEN_669 = inputAdvance ? inputMemBlock_156 : _GEN_156;
  assign _GEN_670 = inputAdvance ? inputMemBlock_157 : _GEN_157;
  assign _GEN_671 = inputAdvance ? inputMemBlock_158 : _GEN_158;
  assign _GEN_672 = inputAdvance ? inputMemBlock_159 : _GEN_159;
  assign _GEN_673 = inputAdvance ? inputMemBlock_160 : _GEN_160;
  assign _GEN_674 = inputAdvance ? inputMemBlock_161 : _GEN_161;
  assign _GEN_675 = inputAdvance ? inputMemBlock_162 : _GEN_162;
  assign _GEN_676 = inputAdvance ? inputMemBlock_163 : _GEN_163;
  assign _GEN_677 = inputAdvance ? inputMemBlock_164 : _GEN_164;
  assign _GEN_678 = inputAdvance ? inputMemBlock_165 : _GEN_165;
  assign _GEN_679 = inputAdvance ? inputMemBlock_166 : _GEN_166;
  assign _GEN_680 = inputAdvance ? inputMemBlock_167 : _GEN_167;
  assign _GEN_681 = inputAdvance ? inputMemBlock_168 : _GEN_168;
  assign _GEN_682 = inputAdvance ? inputMemBlock_169 : _GEN_169;
  assign _GEN_683 = inputAdvance ? inputMemBlock_170 : _GEN_170;
  assign _GEN_684 = inputAdvance ? inputMemBlock_171 : _GEN_171;
  assign _GEN_685 = inputAdvance ? inputMemBlock_172 : _GEN_172;
  assign _GEN_686 = inputAdvance ? inputMemBlock_173 : _GEN_173;
  assign _GEN_687 = inputAdvance ? inputMemBlock_174 : _GEN_174;
  assign _GEN_688 = inputAdvance ? inputMemBlock_175 : _GEN_175;
  assign _GEN_689 = inputAdvance ? inputMemBlock_176 : _GEN_176;
  assign _GEN_690 = inputAdvance ? inputMemBlock_177 : _GEN_177;
  assign _GEN_691 = inputAdvance ? inputMemBlock_178 : _GEN_178;
  assign _GEN_692 = inputAdvance ? inputMemBlock_179 : _GEN_179;
  assign _GEN_693 = inputAdvance ? inputMemBlock_180 : _GEN_180;
  assign _GEN_694 = inputAdvance ? inputMemBlock_181 : _GEN_181;
  assign _GEN_695 = inputAdvance ? inputMemBlock_182 : _GEN_182;
  assign _GEN_696 = inputAdvance ? inputMemBlock_183 : _GEN_183;
  assign _GEN_697 = inputAdvance ? inputMemBlock_184 : _GEN_184;
  assign _GEN_698 = inputAdvance ? inputMemBlock_185 : _GEN_185;
  assign _GEN_699 = inputAdvance ? inputMemBlock_186 : _GEN_186;
  assign _GEN_700 = inputAdvance ? inputMemBlock_187 : _GEN_187;
  assign _GEN_701 = inputAdvance ? inputMemBlock_188 : _GEN_188;
  assign _GEN_702 = inputAdvance ? inputMemBlock_189 : _GEN_189;
  assign _GEN_703 = inputAdvance ? inputMemBlock_190 : _GEN_190;
  assign _GEN_704 = inputAdvance ? inputMemBlock_191 : _GEN_191;
  assign _GEN_705 = inputAdvance ? inputMemBlock_192 : _GEN_192;
  assign _GEN_706 = inputAdvance ? inputMemBlock_193 : _GEN_193;
  assign _GEN_707 = inputAdvance ? inputMemBlock_194 : _GEN_194;
  assign _GEN_708 = inputAdvance ? inputMemBlock_195 : _GEN_195;
  assign _GEN_709 = inputAdvance ? inputMemBlock_196 : _GEN_196;
  assign _GEN_710 = inputAdvance ? inputMemBlock_197 : _GEN_197;
  assign _GEN_711 = inputAdvance ? inputMemBlock_198 : _GEN_198;
  assign _GEN_712 = inputAdvance ? inputMemBlock_199 : _GEN_199;
  assign _GEN_713 = inputAdvance ? inputMemBlock_200 : _GEN_200;
  assign _GEN_714 = inputAdvance ? inputMemBlock_201 : _GEN_201;
  assign _GEN_715 = inputAdvance ? inputMemBlock_202 : _GEN_202;
  assign _GEN_716 = inputAdvance ? inputMemBlock_203 : _GEN_203;
  assign _GEN_717 = inputAdvance ? inputMemBlock_204 : _GEN_204;
  assign _GEN_718 = inputAdvance ? inputMemBlock_205 : _GEN_205;
  assign _GEN_719 = inputAdvance ? inputMemBlock_206 : _GEN_206;
  assign _GEN_720 = inputAdvance ? inputMemBlock_207 : _GEN_207;
  assign _GEN_721 = inputAdvance ? inputMemBlock_208 : _GEN_208;
  assign _GEN_722 = inputAdvance ? inputMemBlock_209 : _GEN_209;
  assign _GEN_723 = inputAdvance ? inputMemBlock_210 : _GEN_210;
  assign _GEN_724 = inputAdvance ? inputMemBlock_211 : _GEN_211;
  assign _GEN_725 = inputAdvance ? inputMemBlock_212 : _GEN_212;
  assign _GEN_726 = inputAdvance ? inputMemBlock_213 : _GEN_213;
  assign _GEN_727 = inputAdvance ? inputMemBlock_214 : _GEN_214;
  assign _GEN_728 = inputAdvance ? inputMemBlock_215 : _GEN_215;
  assign _GEN_729 = inputAdvance ? inputMemBlock_216 : _GEN_216;
  assign _GEN_730 = inputAdvance ? inputMemBlock_217 : _GEN_217;
  assign _GEN_731 = inputAdvance ? inputMemBlock_218 : _GEN_218;
  assign _GEN_732 = inputAdvance ? inputMemBlock_219 : _GEN_219;
  assign _GEN_733 = inputAdvance ? inputMemBlock_220 : _GEN_220;
  assign _GEN_734 = inputAdvance ? inputMemBlock_221 : _GEN_221;
  assign _GEN_735 = inputAdvance ? inputMemBlock_222 : _GEN_222;
  assign _GEN_736 = inputAdvance ? inputMemBlock_223 : _GEN_223;
  assign _GEN_737 = inputAdvance ? inputMemBlock_224 : _GEN_224;
  assign _GEN_738 = inputAdvance ? inputMemBlock_225 : _GEN_225;
  assign _GEN_739 = inputAdvance ? inputMemBlock_226 : _GEN_226;
  assign _GEN_740 = inputAdvance ? inputMemBlock_227 : _GEN_227;
  assign _GEN_741 = inputAdvance ? inputMemBlock_228 : _GEN_228;
  assign _GEN_742 = inputAdvance ? inputMemBlock_229 : _GEN_229;
  assign _GEN_743 = inputAdvance ? inputMemBlock_230 : _GEN_230;
  assign _GEN_744 = inputAdvance ? inputMemBlock_231 : _GEN_231;
  assign _GEN_745 = inputAdvance ? inputMemBlock_232 : _GEN_232;
  assign _GEN_746 = inputAdvance ? inputMemBlock_233 : _GEN_233;
  assign _GEN_747 = inputAdvance ? inputMemBlock_234 : _GEN_234;
  assign _GEN_748 = inputAdvance ? inputMemBlock_235 : _GEN_235;
  assign _GEN_749 = inputAdvance ? inputMemBlock_236 : _GEN_236;
  assign _GEN_750 = inputAdvance ? inputMemBlock_237 : _GEN_237;
  assign _GEN_751 = inputAdvance ? inputMemBlock_238 : _GEN_238;
  assign _GEN_752 = inputAdvance ? inputMemBlock_239 : _GEN_239;
  assign _GEN_753 = inputAdvance ? inputMemBlock_240 : _GEN_240;
  assign _GEN_754 = inputAdvance ? inputMemBlock_241 : _GEN_241;
  assign _GEN_755 = inputAdvance ? inputMemBlock_242 : _GEN_242;
  assign _GEN_756 = inputAdvance ? inputMemBlock_243 : _GEN_243;
  assign _GEN_757 = inputAdvance ? inputMemBlock_244 : _GEN_244;
  assign _GEN_758 = inputAdvance ? inputMemBlock_245 : _GEN_245;
  assign _GEN_759 = inputAdvance ? inputMemBlock_246 : _GEN_246;
  assign _GEN_760 = inputAdvance ? inputMemBlock_247 : _GEN_247;
  assign _GEN_761 = inputAdvance ? inputMemBlock_248 : _GEN_248;
  assign _GEN_762 = inputAdvance ? inputMemBlock_249 : _GEN_249;
  assign _GEN_763 = inputAdvance ? inputMemBlock_250 : _GEN_250;
  assign _GEN_764 = inputAdvance ? inputMemBlock_251 : _GEN_251;
  assign _GEN_765 = inputAdvance ? inputMemBlock_252 : _GEN_252;
  assign _GEN_766 = inputAdvance ? inputMemBlock_253 : _GEN_253;
  assign _GEN_767 = inputAdvance ? inputMemBlock_254 : _GEN_254;
  assign _GEN_768 = inputAdvance ? inputMemBlock_255 : _GEN_255;
  assign _GEN_769 = inputAdvance ? inputMemBlock_256 : _GEN_256;
  assign _GEN_770 = inputAdvance ? inputMemBlock_257 : _GEN_257;
  assign _GEN_771 = inputAdvance ? inputMemBlock_258 : _GEN_258;
  assign _GEN_772 = inputAdvance ? inputMemBlock_259 : _GEN_259;
  assign _GEN_773 = inputAdvance ? inputMemBlock_260 : _GEN_260;
  assign _GEN_774 = inputAdvance ? inputMemBlock_261 : _GEN_261;
  assign _GEN_775 = inputAdvance ? inputMemBlock_262 : _GEN_262;
  assign _GEN_776 = inputAdvance ? inputMemBlock_263 : _GEN_263;
  assign _GEN_777 = inputAdvance ? inputMemBlock_264 : _GEN_264;
  assign _GEN_778 = inputAdvance ? inputMemBlock_265 : _GEN_265;
  assign _GEN_779 = inputAdvance ? inputMemBlock_266 : _GEN_266;
  assign _GEN_780 = inputAdvance ? inputMemBlock_267 : _GEN_267;
  assign _GEN_781 = inputAdvance ? inputMemBlock_268 : _GEN_268;
  assign _GEN_782 = inputAdvance ? inputMemBlock_269 : _GEN_269;
  assign _GEN_783 = inputAdvance ? inputMemBlock_270 : _GEN_270;
  assign _GEN_784 = inputAdvance ? inputMemBlock_271 : _GEN_271;
  assign _GEN_785 = inputAdvance ? inputMemBlock_272 : _GEN_272;
  assign _GEN_786 = inputAdvance ? inputMemBlock_273 : _GEN_273;
  assign _GEN_787 = inputAdvance ? inputMemBlock_274 : _GEN_274;
  assign _GEN_788 = inputAdvance ? inputMemBlock_275 : _GEN_275;
  assign _GEN_789 = inputAdvance ? inputMemBlock_276 : _GEN_276;
  assign _GEN_790 = inputAdvance ? inputMemBlock_277 : _GEN_277;
  assign _GEN_791 = inputAdvance ? inputMemBlock_278 : _GEN_278;
  assign _GEN_792 = inputAdvance ? inputMemBlock_279 : _GEN_279;
  assign _GEN_793 = inputAdvance ? inputMemBlock_280 : _GEN_280;
  assign _GEN_794 = inputAdvance ? inputMemBlock_281 : _GEN_281;
  assign _GEN_795 = inputAdvance ? inputMemBlock_282 : _GEN_282;
  assign _GEN_796 = inputAdvance ? inputMemBlock_283 : _GEN_283;
  assign _GEN_797 = inputAdvance ? inputMemBlock_284 : _GEN_284;
  assign _GEN_798 = inputAdvance ? inputMemBlock_285 : _GEN_285;
  assign _GEN_799 = inputAdvance ? inputMemBlock_286 : _GEN_286;
  assign _GEN_800 = inputAdvance ? inputMemBlock_287 : _GEN_287;
  assign _GEN_801 = inputAdvance ? inputMemBlock_288 : _GEN_288;
  assign _GEN_802 = inputAdvance ? inputMemBlock_289 : _GEN_289;
  assign _GEN_803 = inputAdvance ? inputMemBlock_290 : _GEN_290;
  assign _GEN_804 = inputAdvance ? inputMemBlock_291 : _GEN_291;
  assign _GEN_805 = inputAdvance ? inputMemBlock_292 : _GEN_292;
  assign _GEN_806 = inputAdvance ? inputMemBlock_293 : _GEN_293;
  assign _GEN_807 = inputAdvance ? inputMemBlock_294 : _GEN_294;
  assign _GEN_808 = inputAdvance ? inputMemBlock_295 : _GEN_295;
  assign _GEN_809 = inputAdvance ? inputMemBlock_296 : _GEN_296;
  assign _GEN_810 = inputAdvance ? inputMemBlock_297 : _GEN_297;
  assign _GEN_811 = inputAdvance ? inputMemBlock_298 : _GEN_298;
  assign _GEN_812 = inputAdvance ? inputMemBlock_299 : _GEN_299;
  assign _GEN_813 = inputAdvance ? inputMemBlock_300 : _GEN_300;
  assign _GEN_814 = inputAdvance ? inputMemBlock_301 : _GEN_301;
  assign _GEN_815 = inputAdvance ? inputMemBlock_302 : _GEN_302;
  assign _GEN_816 = inputAdvance ? inputMemBlock_303 : _GEN_303;
  assign _GEN_817 = inputAdvance ? inputMemBlock_304 : _GEN_304;
  assign _GEN_818 = inputAdvance ? inputMemBlock_305 : _GEN_305;
  assign _GEN_819 = inputAdvance ? inputMemBlock_306 : _GEN_306;
  assign _GEN_820 = inputAdvance ? inputMemBlock_307 : _GEN_307;
  assign _GEN_821 = inputAdvance ? inputMemBlock_308 : _GEN_308;
  assign _GEN_822 = inputAdvance ? inputMemBlock_309 : _GEN_309;
  assign _GEN_823 = inputAdvance ? inputMemBlock_310 : _GEN_310;
  assign _GEN_824 = inputAdvance ? inputMemBlock_311 : _GEN_311;
  assign _GEN_825 = inputAdvance ? inputMemBlock_312 : _GEN_312;
  assign _GEN_826 = inputAdvance ? inputMemBlock_313 : _GEN_313;
  assign _GEN_827 = inputAdvance ? inputMemBlock_314 : _GEN_314;
  assign _GEN_828 = inputAdvance ? inputMemBlock_315 : _GEN_315;
  assign _GEN_829 = inputAdvance ? inputMemBlock_316 : _GEN_316;
  assign _GEN_830 = inputAdvance ? inputMemBlock_317 : _GEN_317;
  assign _GEN_831 = inputAdvance ? inputMemBlock_318 : _GEN_318;
  assign _GEN_832 = inputAdvance ? inputMemBlock_319 : _GEN_319;
  assign _GEN_833 = inputAdvance ? inputMemBlock_320 : _GEN_320;
  assign _GEN_834 = inputAdvance ? inputMemBlock_321 : _GEN_321;
  assign _GEN_835 = inputAdvance ? inputMemBlock_322 : _GEN_322;
  assign _GEN_836 = inputAdvance ? inputMemBlock_323 : _GEN_323;
  assign _GEN_837 = inputAdvance ? inputMemBlock_324 : _GEN_324;
  assign _GEN_838 = inputAdvance ? inputMemBlock_325 : _GEN_325;
  assign _GEN_839 = inputAdvance ? inputMemBlock_326 : _GEN_326;
  assign _GEN_840 = inputAdvance ? inputMemBlock_327 : _GEN_327;
  assign _GEN_841 = inputAdvance ? inputMemBlock_328 : _GEN_328;
  assign _GEN_842 = inputAdvance ? inputMemBlock_329 : _GEN_329;
  assign _GEN_843 = inputAdvance ? inputMemBlock_330 : _GEN_330;
  assign _GEN_844 = inputAdvance ? inputMemBlock_331 : _GEN_331;
  assign _GEN_845 = inputAdvance ? inputMemBlock_332 : _GEN_332;
  assign _GEN_846 = inputAdvance ? inputMemBlock_333 : _GEN_333;
  assign _GEN_847 = inputAdvance ? inputMemBlock_334 : _GEN_334;
  assign _GEN_848 = inputAdvance ? inputMemBlock_335 : _GEN_335;
  assign _GEN_849 = inputAdvance ? inputMemBlock_336 : _GEN_336;
  assign _GEN_850 = inputAdvance ? inputMemBlock_337 : _GEN_337;
  assign _GEN_851 = inputAdvance ? inputMemBlock_338 : _GEN_338;
  assign _GEN_852 = inputAdvance ? inputMemBlock_339 : _GEN_339;
  assign _GEN_853 = inputAdvance ? inputMemBlock_340 : _GEN_340;
  assign _GEN_854 = inputAdvance ? inputMemBlock_341 : _GEN_341;
  assign _GEN_855 = inputAdvance ? inputMemBlock_342 : _GEN_342;
  assign _GEN_856 = inputAdvance ? inputMemBlock_343 : _GEN_343;
  assign _GEN_857 = inputAdvance ? inputMemBlock_344 : _GEN_344;
  assign _GEN_858 = inputAdvance ? inputMemBlock_345 : _GEN_345;
  assign _GEN_859 = inputAdvance ? inputMemBlock_346 : _GEN_346;
  assign _GEN_860 = inputAdvance ? inputMemBlock_347 : _GEN_347;
  assign _GEN_861 = inputAdvance ? inputMemBlock_348 : _GEN_348;
  assign _GEN_862 = inputAdvance ? inputMemBlock_349 : _GEN_349;
  assign _GEN_863 = inputAdvance ? inputMemBlock_350 : _GEN_350;
  assign _GEN_864 = inputAdvance ? inputMemBlock_351 : _GEN_351;
  assign _GEN_865 = inputAdvance ? inputMemBlock_352 : _GEN_352;
  assign _GEN_866 = inputAdvance ? inputMemBlock_353 : _GEN_353;
  assign _GEN_867 = inputAdvance ? inputMemBlock_354 : _GEN_354;
  assign _GEN_868 = inputAdvance ? inputMemBlock_355 : _GEN_355;
  assign _GEN_869 = inputAdvance ? inputMemBlock_356 : _GEN_356;
  assign _GEN_870 = inputAdvance ? inputMemBlock_357 : _GEN_357;
  assign _GEN_871 = inputAdvance ? inputMemBlock_358 : _GEN_358;
  assign _GEN_872 = inputAdvance ? inputMemBlock_359 : _GEN_359;
  assign _GEN_873 = inputAdvance ? inputMemBlock_360 : _GEN_360;
  assign _GEN_874 = inputAdvance ? inputMemBlock_361 : _GEN_361;
  assign _GEN_875 = inputAdvance ? inputMemBlock_362 : _GEN_362;
  assign _GEN_876 = inputAdvance ? inputMemBlock_363 : _GEN_363;
  assign _GEN_877 = inputAdvance ? inputMemBlock_364 : _GEN_364;
  assign _GEN_878 = inputAdvance ? inputMemBlock_365 : _GEN_365;
  assign _GEN_879 = inputAdvance ? inputMemBlock_366 : _GEN_366;
  assign _GEN_880 = inputAdvance ? inputMemBlock_367 : _GEN_367;
  assign _GEN_881 = inputAdvance ? inputMemBlock_368 : _GEN_368;
  assign _GEN_882 = inputAdvance ? inputMemBlock_369 : _GEN_369;
  assign _GEN_883 = inputAdvance ? inputMemBlock_370 : _GEN_370;
  assign _GEN_884 = inputAdvance ? inputMemBlock_371 : _GEN_371;
  assign _GEN_885 = inputAdvance ? inputMemBlock_372 : _GEN_372;
  assign _GEN_886 = inputAdvance ? inputMemBlock_373 : _GEN_373;
  assign _GEN_887 = inputAdvance ? inputMemBlock_374 : _GEN_374;
  assign _GEN_888 = inputAdvance ? inputMemBlock_375 : _GEN_375;
  assign _GEN_889 = inputAdvance ? inputMemBlock_376 : _GEN_376;
  assign _GEN_890 = inputAdvance ? inputMemBlock_377 : _GEN_377;
  assign _GEN_891 = inputAdvance ? inputMemBlock_378 : _GEN_378;
  assign _GEN_892 = inputAdvance ? inputMemBlock_379 : _GEN_379;
  assign _GEN_893 = inputAdvance ? inputMemBlock_380 : _GEN_380;
  assign _GEN_894 = inputAdvance ? inputMemBlock_381 : _GEN_381;
  assign _GEN_895 = inputAdvance ? inputMemBlock_382 : _GEN_382;
  assign _GEN_896 = inputAdvance ? inputMemBlock_383 : _GEN_383;
  assign _GEN_897 = inputAdvance ? inputMemBlock_384 : _GEN_384;
  assign _GEN_898 = inputAdvance ? inputMemBlock_385 : _GEN_385;
  assign _GEN_899 = inputAdvance ? inputMemBlock_386 : _GEN_386;
  assign _GEN_900 = inputAdvance ? inputMemBlock_387 : _GEN_387;
  assign _GEN_901 = inputAdvance ? inputMemBlock_388 : _GEN_388;
  assign _GEN_902 = inputAdvance ? inputMemBlock_389 : _GEN_389;
  assign _GEN_903 = inputAdvance ? inputMemBlock_390 : _GEN_390;
  assign _GEN_904 = inputAdvance ? inputMemBlock_391 : _GEN_391;
  assign _GEN_905 = inputAdvance ? inputMemBlock_392 : _GEN_392;
  assign _GEN_906 = inputAdvance ? inputMemBlock_393 : _GEN_393;
  assign _GEN_907 = inputAdvance ? inputMemBlock_394 : _GEN_394;
  assign _GEN_908 = inputAdvance ? inputMemBlock_395 : _GEN_395;
  assign _GEN_909 = inputAdvance ? inputMemBlock_396 : _GEN_396;
  assign _GEN_910 = inputAdvance ? inputMemBlock_397 : _GEN_397;
  assign _GEN_911 = inputAdvance ? inputMemBlock_398 : _GEN_398;
  assign _GEN_912 = inputAdvance ? inputMemBlock_399 : _GEN_399;
  assign _GEN_913 = inputAdvance ? inputMemBlock_400 : _GEN_400;
  assign _GEN_914 = inputAdvance ? inputMemBlock_401 : _GEN_401;
  assign _GEN_915 = inputAdvance ? inputMemBlock_402 : _GEN_402;
  assign _GEN_916 = inputAdvance ? inputMemBlock_403 : _GEN_403;
  assign _GEN_917 = inputAdvance ? inputMemBlock_404 : _GEN_404;
  assign _GEN_918 = inputAdvance ? inputMemBlock_405 : _GEN_405;
  assign _GEN_919 = inputAdvance ? inputMemBlock_406 : _GEN_406;
  assign _GEN_920 = inputAdvance ? inputMemBlock_407 : _GEN_407;
  assign _GEN_921 = inputAdvance ? inputMemBlock_408 : _GEN_408;
  assign _GEN_922 = inputAdvance ? inputMemBlock_409 : _GEN_409;
  assign _GEN_923 = inputAdvance ? inputMemBlock_410 : _GEN_410;
  assign _GEN_924 = inputAdvance ? inputMemBlock_411 : _GEN_411;
  assign _GEN_925 = inputAdvance ? inputMemBlock_412 : _GEN_412;
  assign _GEN_926 = inputAdvance ? inputMemBlock_413 : _GEN_413;
  assign _GEN_927 = inputAdvance ? inputMemBlock_414 : _GEN_414;
  assign _GEN_928 = inputAdvance ? inputMemBlock_415 : _GEN_415;
  assign _GEN_929 = inputAdvance ? inputMemBlock_416 : _GEN_416;
  assign _GEN_930 = inputAdvance ? inputMemBlock_417 : _GEN_417;
  assign _GEN_931 = inputAdvance ? inputMemBlock_418 : _GEN_418;
  assign _GEN_932 = inputAdvance ? inputMemBlock_419 : _GEN_419;
  assign _GEN_933 = inputAdvance ? inputMemBlock_420 : _GEN_420;
  assign _GEN_934 = inputAdvance ? inputMemBlock_421 : _GEN_421;
  assign _GEN_935 = inputAdvance ? inputMemBlock_422 : _GEN_422;
  assign _GEN_936 = inputAdvance ? inputMemBlock_423 : _GEN_423;
  assign _GEN_937 = inputAdvance ? inputMemBlock_424 : _GEN_424;
  assign _GEN_938 = inputAdvance ? inputMemBlock_425 : _GEN_425;
  assign _GEN_939 = inputAdvance ? inputMemBlock_426 : _GEN_426;
  assign _GEN_940 = inputAdvance ? inputMemBlock_427 : _GEN_427;
  assign _GEN_941 = inputAdvance ? inputMemBlock_428 : _GEN_428;
  assign _GEN_942 = inputAdvance ? inputMemBlock_429 : _GEN_429;
  assign _GEN_943 = inputAdvance ? inputMemBlock_430 : _GEN_430;
  assign _GEN_944 = inputAdvance ? inputMemBlock_431 : _GEN_431;
  assign _GEN_945 = inputAdvance ? inputMemBlock_432 : _GEN_432;
  assign _GEN_946 = inputAdvance ? inputMemBlock_433 : _GEN_433;
  assign _GEN_947 = inputAdvance ? inputMemBlock_434 : _GEN_434;
  assign _GEN_948 = inputAdvance ? inputMemBlock_435 : _GEN_435;
  assign _GEN_949 = inputAdvance ? inputMemBlock_436 : _GEN_436;
  assign _GEN_950 = inputAdvance ? inputMemBlock_437 : _GEN_437;
  assign _GEN_951 = inputAdvance ? inputMemBlock_438 : _GEN_438;
  assign _GEN_952 = inputAdvance ? inputMemBlock_439 : _GEN_439;
  assign _GEN_953 = inputAdvance ? inputMemBlock_440 : _GEN_440;
  assign _GEN_954 = inputAdvance ? inputMemBlock_441 : _GEN_441;
  assign _GEN_955 = inputAdvance ? inputMemBlock_442 : _GEN_442;
  assign _GEN_956 = inputAdvance ? inputMemBlock_443 : _GEN_443;
  assign _GEN_957 = inputAdvance ? inputMemBlock_444 : _GEN_444;
  assign _GEN_958 = inputAdvance ? inputMemBlock_445 : _GEN_445;
  assign _GEN_959 = inputAdvance ? inputMemBlock_446 : _GEN_446;
  assign _GEN_960 = inputAdvance ? inputMemBlock_447 : _GEN_447;
  assign _GEN_961 = inputAdvance ? inputMemBlock_448 : _GEN_448;
  assign _GEN_962 = inputAdvance ? inputMemBlock_449 : _GEN_449;
  assign _GEN_963 = inputAdvance ? inputMemBlock_450 : _GEN_450;
  assign _GEN_964 = inputAdvance ? inputMemBlock_451 : _GEN_451;
  assign _GEN_965 = inputAdvance ? inputMemBlock_452 : _GEN_452;
  assign _GEN_966 = inputAdvance ? inputMemBlock_453 : _GEN_453;
  assign _GEN_967 = inputAdvance ? inputMemBlock_454 : _GEN_454;
  assign _GEN_968 = inputAdvance ? inputMemBlock_455 : _GEN_455;
  assign _GEN_969 = inputAdvance ? inputMemBlock_456 : _GEN_456;
  assign _GEN_970 = inputAdvance ? inputMemBlock_457 : _GEN_457;
  assign _GEN_971 = inputAdvance ? inputMemBlock_458 : _GEN_458;
  assign _GEN_972 = inputAdvance ? inputMemBlock_459 : _GEN_459;
  assign _GEN_973 = inputAdvance ? inputMemBlock_460 : _GEN_460;
  assign _GEN_974 = inputAdvance ? inputMemBlock_461 : _GEN_461;
  assign _GEN_975 = inputAdvance ? inputMemBlock_462 : _GEN_462;
  assign _GEN_976 = inputAdvance ? inputMemBlock_463 : _GEN_463;
  assign _GEN_977 = inputAdvance ? inputMemBlock_464 : _GEN_464;
  assign _GEN_978 = inputAdvance ? inputMemBlock_465 : _GEN_465;
  assign _GEN_979 = inputAdvance ? inputMemBlock_466 : _GEN_466;
  assign _GEN_980 = inputAdvance ? inputMemBlock_467 : _GEN_467;
  assign _GEN_981 = inputAdvance ? inputMemBlock_468 : _GEN_468;
  assign _GEN_982 = inputAdvance ? inputMemBlock_469 : _GEN_469;
  assign _GEN_983 = inputAdvance ? inputMemBlock_470 : _GEN_470;
  assign _GEN_984 = inputAdvance ? inputMemBlock_471 : _GEN_471;
  assign _GEN_985 = inputAdvance ? inputMemBlock_472 : _GEN_472;
  assign _GEN_986 = inputAdvance ? inputMemBlock_473 : _GEN_473;
  assign _GEN_987 = inputAdvance ? inputMemBlock_474 : _GEN_474;
  assign _GEN_988 = inputAdvance ? inputMemBlock_475 : _GEN_475;
  assign _GEN_989 = inputAdvance ? inputMemBlock_476 : _GEN_476;
  assign _GEN_990 = inputAdvance ? inputMemBlock_477 : _GEN_477;
  assign _GEN_991 = inputAdvance ? inputMemBlock_478 : _GEN_478;
  assign _GEN_992 = inputAdvance ? inputMemBlock_479 : _GEN_479;
  assign _GEN_993 = inputAdvance ? inputMemBlock_480 : _GEN_480;
  assign _GEN_994 = inputAdvance ? inputMemBlock_481 : _GEN_481;
  assign _GEN_995 = inputAdvance ? inputMemBlock_482 : _GEN_482;
  assign _GEN_996 = inputAdvance ? inputMemBlock_483 : _GEN_483;
  assign _GEN_997 = inputAdvance ? inputMemBlock_484 : _GEN_484;
  assign _GEN_998 = inputAdvance ? inputMemBlock_485 : _GEN_485;
  assign _GEN_999 = inputAdvance ? inputMemBlock_486 : _GEN_486;
  assign _GEN_1000 = inputAdvance ? inputMemBlock_487 : _GEN_487;
  assign _GEN_1001 = inputAdvance ? inputMemBlock_488 : _GEN_488;
  assign _GEN_1002 = inputAdvance ? inputMemBlock_489 : _GEN_489;
  assign _GEN_1003 = inputAdvance ? inputMemBlock_490 : _GEN_490;
  assign _GEN_1004 = inputAdvance ? inputMemBlock_491 : _GEN_491;
  assign _GEN_1005 = inputAdvance ? inputMemBlock_492 : _GEN_492;
  assign _GEN_1006 = inputAdvance ? inputMemBlock_493 : _GEN_493;
  assign _GEN_1007 = inputAdvance ? inputMemBlock_494 : _GEN_494;
  assign _GEN_1008 = inputAdvance ? inputMemBlock_495 : _GEN_495;
  assign _GEN_1009 = inputAdvance ? inputMemBlock_496 : _GEN_496;
  assign _GEN_1010 = inputAdvance ? inputMemBlock_497 : _GEN_497;
  assign _GEN_1011 = inputAdvance ? inputMemBlock_498 : _GEN_498;
  assign _GEN_1012 = inputAdvance ? inputMemBlock_499 : _GEN_499;
  assign _GEN_1013 = inputAdvance ? inputMemBlock_500 : _GEN_500;
  assign _GEN_1014 = inputAdvance ? inputMemBlock_501 : _GEN_501;
  assign _GEN_1015 = inputAdvance ? inputMemBlock_502 : _GEN_502;
  assign _GEN_1016 = inputAdvance ? inputMemBlock_503 : _GEN_503;
  assign _GEN_1017 = inputAdvance ? inputMemBlock_504 : _GEN_504;
  assign _GEN_1018 = inputAdvance ? inputMemBlock_505 : _GEN_505;
  assign _GEN_1019 = inputAdvance ? inputMemBlock_506 : _GEN_506;
  assign _GEN_1020 = inputAdvance ? inputMemBlock_507 : _GEN_507;
  assign _GEN_1021 = inputAdvance ? inputMemBlock_508 : _GEN_508;
  assign _GEN_1022 = inputAdvance ? inputMemBlock_509 : _GEN_509;
  assign _GEN_1023 = inputAdvance ? inputMemBlock_510 : _GEN_510;
  assign _GEN_1024 = inputAdvance ? inputMemBlock_511 : _GEN_511;
  assign _T_1587 = outputBits + 10'h1;
  assign _T_1588 = _T_1587[9:0];
  assign _GEN_1025 = nextBitValid ? nextBit : outputMemBlock_511;
  assign _GEN_1026 = nextBitValid ? outputMemBlock_1 : outputMemBlock_0;
  assign _GEN_1027 = nextBitValid ? outputMemBlock_2 : outputMemBlock_1;
  assign _GEN_1028 = nextBitValid ? outputMemBlock_3 : outputMemBlock_2;
  assign _GEN_1029 = nextBitValid ? outputMemBlock_4 : outputMemBlock_3;
  assign _GEN_1030 = nextBitValid ? outputMemBlock_5 : outputMemBlock_4;
  assign _GEN_1031 = nextBitValid ? outputMemBlock_6 : outputMemBlock_5;
  assign _GEN_1032 = nextBitValid ? outputMemBlock_7 : outputMemBlock_6;
  assign _GEN_1033 = nextBitValid ? outputMemBlock_8 : outputMemBlock_7;
  assign _GEN_1034 = nextBitValid ? outputMemBlock_9 : outputMemBlock_8;
  assign _GEN_1035 = nextBitValid ? outputMemBlock_10 : outputMemBlock_9;
  assign _GEN_1036 = nextBitValid ? outputMemBlock_11 : outputMemBlock_10;
  assign _GEN_1037 = nextBitValid ? outputMemBlock_12 : outputMemBlock_11;
  assign _GEN_1038 = nextBitValid ? outputMemBlock_13 : outputMemBlock_12;
  assign _GEN_1039 = nextBitValid ? outputMemBlock_14 : outputMemBlock_13;
  assign _GEN_1040 = nextBitValid ? outputMemBlock_15 : outputMemBlock_14;
  assign _GEN_1041 = nextBitValid ? outputMemBlock_16 : outputMemBlock_15;
  assign _GEN_1042 = nextBitValid ? outputMemBlock_17 : outputMemBlock_16;
  assign _GEN_1043 = nextBitValid ? outputMemBlock_18 : outputMemBlock_17;
  assign _GEN_1044 = nextBitValid ? outputMemBlock_19 : outputMemBlock_18;
  assign _GEN_1045 = nextBitValid ? outputMemBlock_20 : outputMemBlock_19;
  assign _GEN_1046 = nextBitValid ? outputMemBlock_21 : outputMemBlock_20;
  assign _GEN_1047 = nextBitValid ? outputMemBlock_22 : outputMemBlock_21;
  assign _GEN_1048 = nextBitValid ? outputMemBlock_23 : outputMemBlock_22;
  assign _GEN_1049 = nextBitValid ? outputMemBlock_24 : outputMemBlock_23;
  assign _GEN_1050 = nextBitValid ? outputMemBlock_25 : outputMemBlock_24;
  assign _GEN_1051 = nextBitValid ? outputMemBlock_26 : outputMemBlock_25;
  assign _GEN_1052 = nextBitValid ? outputMemBlock_27 : outputMemBlock_26;
  assign _GEN_1053 = nextBitValid ? outputMemBlock_28 : outputMemBlock_27;
  assign _GEN_1054 = nextBitValid ? outputMemBlock_29 : outputMemBlock_28;
  assign _GEN_1055 = nextBitValid ? outputMemBlock_30 : outputMemBlock_29;
  assign _GEN_1056 = nextBitValid ? outputMemBlock_31 : outputMemBlock_30;
  assign _GEN_1057 = nextBitValid ? outputMemBlock_32 : outputMemBlock_31;
  assign _GEN_1058 = nextBitValid ? outputMemBlock_33 : outputMemBlock_32;
  assign _GEN_1059 = nextBitValid ? outputMemBlock_34 : outputMemBlock_33;
  assign _GEN_1060 = nextBitValid ? outputMemBlock_35 : outputMemBlock_34;
  assign _GEN_1061 = nextBitValid ? outputMemBlock_36 : outputMemBlock_35;
  assign _GEN_1062 = nextBitValid ? outputMemBlock_37 : outputMemBlock_36;
  assign _GEN_1063 = nextBitValid ? outputMemBlock_38 : outputMemBlock_37;
  assign _GEN_1064 = nextBitValid ? outputMemBlock_39 : outputMemBlock_38;
  assign _GEN_1065 = nextBitValid ? outputMemBlock_40 : outputMemBlock_39;
  assign _GEN_1066 = nextBitValid ? outputMemBlock_41 : outputMemBlock_40;
  assign _GEN_1067 = nextBitValid ? outputMemBlock_42 : outputMemBlock_41;
  assign _GEN_1068 = nextBitValid ? outputMemBlock_43 : outputMemBlock_42;
  assign _GEN_1069 = nextBitValid ? outputMemBlock_44 : outputMemBlock_43;
  assign _GEN_1070 = nextBitValid ? outputMemBlock_45 : outputMemBlock_44;
  assign _GEN_1071 = nextBitValid ? outputMemBlock_46 : outputMemBlock_45;
  assign _GEN_1072 = nextBitValid ? outputMemBlock_47 : outputMemBlock_46;
  assign _GEN_1073 = nextBitValid ? outputMemBlock_48 : outputMemBlock_47;
  assign _GEN_1074 = nextBitValid ? outputMemBlock_49 : outputMemBlock_48;
  assign _GEN_1075 = nextBitValid ? outputMemBlock_50 : outputMemBlock_49;
  assign _GEN_1076 = nextBitValid ? outputMemBlock_51 : outputMemBlock_50;
  assign _GEN_1077 = nextBitValid ? outputMemBlock_52 : outputMemBlock_51;
  assign _GEN_1078 = nextBitValid ? outputMemBlock_53 : outputMemBlock_52;
  assign _GEN_1079 = nextBitValid ? outputMemBlock_54 : outputMemBlock_53;
  assign _GEN_1080 = nextBitValid ? outputMemBlock_55 : outputMemBlock_54;
  assign _GEN_1081 = nextBitValid ? outputMemBlock_56 : outputMemBlock_55;
  assign _GEN_1082 = nextBitValid ? outputMemBlock_57 : outputMemBlock_56;
  assign _GEN_1083 = nextBitValid ? outputMemBlock_58 : outputMemBlock_57;
  assign _GEN_1084 = nextBitValid ? outputMemBlock_59 : outputMemBlock_58;
  assign _GEN_1085 = nextBitValid ? outputMemBlock_60 : outputMemBlock_59;
  assign _GEN_1086 = nextBitValid ? outputMemBlock_61 : outputMemBlock_60;
  assign _GEN_1087 = nextBitValid ? outputMemBlock_62 : outputMemBlock_61;
  assign _GEN_1088 = nextBitValid ? outputMemBlock_63 : outputMemBlock_62;
  assign _GEN_1089 = nextBitValid ? outputMemBlock_64 : outputMemBlock_63;
  assign _GEN_1090 = nextBitValid ? outputMemBlock_65 : outputMemBlock_64;
  assign _GEN_1091 = nextBitValid ? outputMemBlock_66 : outputMemBlock_65;
  assign _GEN_1092 = nextBitValid ? outputMemBlock_67 : outputMemBlock_66;
  assign _GEN_1093 = nextBitValid ? outputMemBlock_68 : outputMemBlock_67;
  assign _GEN_1094 = nextBitValid ? outputMemBlock_69 : outputMemBlock_68;
  assign _GEN_1095 = nextBitValid ? outputMemBlock_70 : outputMemBlock_69;
  assign _GEN_1096 = nextBitValid ? outputMemBlock_71 : outputMemBlock_70;
  assign _GEN_1097 = nextBitValid ? outputMemBlock_72 : outputMemBlock_71;
  assign _GEN_1098 = nextBitValid ? outputMemBlock_73 : outputMemBlock_72;
  assign _GEN_1099 = nextBitValid ? outputMemBlock_74 : outputMemBlock_73;
  assign _GEN_1100 = nextBitValid ? outputMemBlock_75 : outputMemBlock_74;
  assign _GEN_1101 = nextBitValid ? outputMemBlock_76 : outputMemBlock_75;
  assign _GEN_1102 = nextBitValid ? outputMemBlock_77 : outputMemBlock_76;
  assign _GEN_1103 = nextBitValid ? outputMemBlock_78 : outputMemBlock_77;
  assign _GEN_1104 = nextBitValid ? outputMemBlock_79 : outputMemBlock_78;
  assign _GEN_1105 = nextBitValid ? outputMemBlock_80 : outputMemBlock_79;
  assign _GEN_1106 = nextBitValid ? outputMemBlock_81 : outputMemBlock_80;
  assign _GEN_1107 = nextBitValid ? outputMemBlock_82 : outputMemBlock_81;
  assign _GEN_1108 = nextBitValid ? outputMemBlock_83 : outputMemBlock_82;
  assign _GEN_1109 = nextBitValid ? outputMemBlock_84 : outputMemBlock_83;
  assign _GEN_1110 = nextBitValid ? outputMemBlock_85 : outputMemBlock_84;
  assign _GEN_1111 = nextBitValid ? outputMemBlock_86 : outputMemBlock_85;
  assign _GEN_1112 = nextBitValid ? outputMemBlock_87 : outputMemBlock_86;
  assign _GEN_1113 = nextBitValid ? outputMemBlock_88 : outputMemBlock_87;
  assign _GEN_1114 = nextBitValid ? outputMemBlock_89 : outputMemBlock_88;
  assign _GEN_1115 = nextBitValid ? outputMemBlock_90 : outputMemBlock_89;
  assign _GEN_1116 = nextBitValid ? outputMemBlock_91 : outputMemBlock_90;
  assign _GEN_1117 = nextBitValid ? outputMemBlock_92 : outputMemBlock_91;
  assign _GEN_1118 = nextBitValid ? outputMemBlock_93 : outputMemBlock_92;
  assign _GEN_1119 = nextBitValid ? outputMemBlock_94 : outputMemBlock_93;
  assign _GEN_1120 = nextBitValid ? outputMemBlock_95 : outputMemBlock_94;
  assign _GEN_1121 = nextBitValid ? outputMemBlock_96 : outputMemBlock_95;
  assign _GEN_1122 = nextBitValid ? outputMemBlock_97 : outputMemBlock_96;
  assign _GEN_1123 = nextBitValid ? outputMemBlock_98 : outputMemBlock_97;
  assign _GEN_1124 = nextBitValid ? outputMemBlock_99 : outputMemBlock_98;
  assign _GEN_1125 = nextBitValid ? outputMemBlock_100 : outputMemBlock_99;
  assign _GEN_1126 = nextBitValid ? outputMemBlock_101 : outputMemBlock_100;
  assign _GEN_1127 = nextBitValid ? outputMemBlock_102 : outputMemBlock_101;
  assign _GEN_1128 = nextBitValid ? outputMemBlock_103 : outputMemBlock_102;
  assign _GEN_1129 = nextBitValid ? outputMemBlock_104 : outputMemBlock_103;
  assign _GEN_1130 = nextBitValid ? outputMemBlock_105 : outputMemBlock_104;
  assign _GEN_1131 = nextBitValid ? outputMemBlock_106 : outputMemBlock_105;
  assign _GEN_1132 = nextBitValid ? outputMemBlock_107 : outputMemBlock_106;
  assign _GEN_1133 = nextBitValid ? outputMemBlock_108 : outputMemBlock_107;
  assign _GEN_1134 = nextBitValid ? outputMemBlock_109 : outputMemBlock_108;
  assign _GEN_1135 = nextBitValid ? outputMemBlock_110 : outputMemBlock_109;
  assign _GEN_1136 = nextBitValid ? outputMemBlock_111 : outputMemBlock_110;
  assign _GEN_1137 = nextBitValid ? outputMemBlock_112 : outputMemBlock_111;
  assign _GEN_1138 = nextBitValid ? outputMemBlock_113 : outputMemBlock_112;
  assign _GEN_1139 = nextBitValid ? outputMemBlock_114 : outputMemBlock_113;
  assign _GEN_1140 = nextBitValid ? outputMemBlock_115 : outputMemBlock_114;
  assign _GEN_1141 = nextBitValid ? outputMemBlock_116 : outputMemBlock_115;
  assign _GEN_1142 = nextBitValid ? outputMemBlock_117 : outputMemBlock_116;
  assign _GEN_1143 = nextBitValid ? outputMemBlock_118 : outputMemBlock_117;
  assign _GEN_1144 = nextBitValid ? outputMemBlock_119 : outputMemBlock_118;
  assign _GEN_1145 = nextBitValid ? outputMemBlock_120 : outputMemBlock_119;
  assign _GEN_1146 = nextBitValid ? outputMemBlock_121 : outputMemBlock_120;
  assign _GEN_1147 = nextBitValid ? outputMemBlock_122 : outputMemBlock_121;
  assign _GEN_1148 = nextBitValid ? outputMemBlock_123 : outputMemBlock_122;
  assign _GEN_1149 = nextBitValid ? outputMemBlock_124 : outputMemBlock_123;
  assign _GEN_1150 = nextBitValid ? outputMemBlock_125 : outputMemBlock_124;
  assign _GEN_1151 = nextBitValid ? outputMemBlock_126 : outputMemBlock_125;
  assign _GEN_1152 = nextBitValid ? outputMemBlock_127 : outputMemBlock_126;
  assign _GEN_1153 = nextBitValid ? outputMemBlock_128 : outputMemBlock_127;
  assign _GEN_1154 = nextBitValid ? outputMemBlock_129 : outputMemBlock_128;
  assign _GEN_1155 = nextBitValid ? outputMemBlock_130 : outputMemBlock_129;
  assign _GEN_1156 = nextBitValid ? outputMemBlock_131 : outputMemBlock_130;
  assign _GEN_1157 = nextBitValid ? outputMemBlock_132 : outputMemBlock_131;
  assign _GEN_1158 = nextBitValid ? outputMemBlock_133 : outputMemBlock_132;
  assign _GEN_1159 = nextBitValid ? outputMemBlock_134 : outputMemBlock_133;
  assign _GEN_1160 = nextBitValid ? outputMemBlock_135 : outputMemBlock_134;
  assign _GEN_1161 = nextBitValid ? outputMemBlock_136 : outputMemBlock_135;
  assign _GEN_1162 = nextBitValid ? outputMemBlock_137 : outputMemBlock_136;
  assign _GEN_1163 = nextBitValid ? outputMemBlock_138 : outputMemBlock_137;
  assign _GEN_1164 = nextBitValid ? outputMemBlock_139 : outputMemBlock_138;
  assign _GEN_1165 = nextBitValid ? outputMemBlock_140 : outputMemBlock_139;
  assign _GEN_1166 = nextBitValid ? outputMemBlock_141 : outputMemBlock_140;
  assign _GEN_1167 = nextBitValid ? outputMemBlock_142 : outputMemBlock_141;
  assign _GEN_1168 = nextBitValid ? outputMemBlock_143 : outputMemBlock_142;
  assign _GEN_1169 = nextBitValid ? outputMemBlock_144 : outputMemBlock_143;
  assign _GEN_1170 = nextBitValid ? outputMemBlock_145 : outputMemBlock_144;
  assign _GEN_1171 = nextBitValid ? outputMemBlock_146 : outputMemBlock_145;
  assign _GEN_1172 = nextBitValid ? outputMemBlock_147 : outputMemBlock_146;
  assign _GEN_1173 = nextBitValid ? outputMemBlock_148 : outputMemBlock_147;
  assign _GEN_1174 = nextBitValid ? outputMemBlock_149 : outputMemBlock_148;
  assign _GEN_1175 = nextBitValid ? outputMemBlock_150 : outputMemBlock_149;
  assign _GEN_1176 = nextBitValid ? outputMemBlock_151 : outputMemBlock_150;
  assign _GEN_1177 = nextBitValid ? outputMemBlock_152 : outputMemBlock_151;
  assign _GEN_1178 = nextBitValid ? outputMemBlock_153 : outputMemBlock_152;
  assign _GEN_1179 = nextBitValid ? outputMemBlock_154 : outputMemBlock_153;
  assign _GEN_1180 = nextBitValid ? outputMemBlock_155 : outputMemBlock_154;
  assign _GEN_1181 = nextBitValid ? outputMemBlock_156 : outputMemBlock_155;
  assign _GEN_1182 = nextBitValid ? outputMemBlock_157 : outputMemBlock_156;
  assign _GEN_1183 = nextBitValid ? outputMemBlock_158 : outputMemBlock_157;
  assign _GEN_1184 = nextBitValid ? outputMemBlock_159 : outputMemBlock_158;
  assign _GEN_1185 = nextBitValid ? outputMemBlock_160 : outputMemBlock_159;
  assign _GEN_1186 = nextBitValid ? outputMemBlock_161 : outputMemBlock_160;
  assign _GEN_1187 = nextBitValid ? outputMemBlock_162 : outputMemBlock_161;
  assign _GEN_1188 = nextBitValid ? outputMemBlock_163 : outputMemBlock_162;
  assign _GEN_1189 = nextBitValid ? outputMemBlock_164 : outputMemBlock_163;
  assign _GEN_1190 = nextBitValid ? outputMemBlock_165 : outputMemBlock_164;
  assign _GEN_1191 = nextBitValid ? outputMemBlock_166 : outputMemBlock_165;
  assign _GEN_1192 = nextBitValid ? outputMemBlock_167 : outputMemBlock_166;
  assign _GEN_1193 = nextBitValid ? outputMemBlock_168 : outputMemBlock_167;
  assign _GEN_1194 = nextBitValid ? outputMemBlock_169 : outputMemBlock_168;
  assign _GEN_1195 = nextBitValid ? outputMemBlock_170 : outputMemBlock_169;
  assign _GEN_1196 = nextBitValid ? outputMemBlock_171 : outputMemBlock_170;
  assign _GEN_1197 = nextBitValid ? outputMemBlock_172 : outputMemBlock_171;
  assign _GEN_1198 = nextBitValid ? outputMemBlock_173 : outputMemBlock_172;
  assign _GEN_1199 = nextBitValid ? outputMemBlock_174 : outputMemBlock_173;
  assign _GEN_1200 = nextBitValid ? outputMemBlock_175 : outputMemBlock_174;
  assign _GEN_1201 = nextBitValid ? outputMemBlock_176 : outputMemBlock_175;
  assign _GEN_1202 = nextBitValid ? outputMemBlock_177 : outputMemBlock_176;
  assign _GEN_1203 = nextBitValid ? outputMemBlock_178 : outputMemBlock_177;
  assign _GEN_1204 = nextBitValid ? outputMemBlock_179 : outputMemBlock_178;
  assign _GEN_1205 = nextBitValid ? outputMemBlock_180 : outputMemBlock_179;
  assign _GEN_1206 = nextBitValid ? outputMemBlock_181 : outputMemBlock_180;
  assign _GEN_1207 = nextBitValid ? outputMemBlock_182 : outputMemBlock_181;
  assign _GEN_1208 = nextBitValid ? outputMemBlock_183 : outputMemBlock_182;
  assign _GEN_1209 = nextBitValid ? outputMemBlock_184 : outputMemBlock_183;
  assign _GEN_1210 = nextBitValid ? outputMemBlock_185 : outputMemBlock_184;
  assign _GEN_1211 = nextBitValid ? outputMemBlock_186 : outputMemBlock_185;
  assign _GEN_1212 = nextBitValid ? outputMemBlock_187 : outputMemBlock_186;
  assign _GEN_1213 = nextBitValid ? outputMemBlock_188 : outputMemBlock_187;
  assign _GEN_1214 = nextBitValid ? outputMemBlock_189 : outputMemBlock_188;
  assign _GEN_1215 = nextBitValid ? outputMemBlock_190 : outputMemBlock_189;
  assign _GEN_1216 = nextBitValid ? outputMemBlock_191 : outputMemBlock_190;
  assign _GEN_1217 = nextBitValid ? outputMemBlock_192 : outputMemBlock_191;
  assign _GEN_1218 = nextBitValid ? outputMemBlock_193 : outputMemBlock_192;
  assign _GEN_1219 = nextBitValid ? outputMemBlock_194 : outputMemBlock_193;
  assign _GEN_1220 = nextBitValid ? outputMemBlock_195 : outputMemBlock_194;
  assign _GEN_1221 = nextBitValid ? outputMemBlock_196 : outputMemBlock_195;
  assign _GEN_1222 = nextBitValid ? outputMemBlock_197 : outputMemBlock_196;
  assign _GEN_1223 = nextBitValid ? outputMemBlock_198 : outputMemBlock_197;
  assign _GEN_1224 = nextBitValid ? outputMemBlock_199 : outputMemBlock_198;
  assign _GEN_1225 = nextBitValid ? outputMemBlock_200 : outputMemBlock_199;
  assign _GEN_1226 = nextBitValid ? outputMemBlock_201 : outputMemBlock_200;
  assign _GEN_1227 = nextBitValid ? outputMemBlock_202 : outputMemBlock_201;
  assign _GEN_1228 = nextBitValid ? outputMemBlock_203 : outputMemBlock_202;
  assign _GEN_1229 = nextBitValid ? outputMemBlock_204 : outputMemBlock_203;
  assign _GEN_1230 = nextBitValid ? outputMemBlock_205 : outputMemBlock_204;
  assign _GEN_1231 = nextBitValid ? outputMemBlock_206 : outputMemBlock_205;
  assign _GEN_1232 = nextBitValid ? outputMemBlock_207 : outputMemBlock_206;
  assign _GEN_1233 = nextBitValid ? outputMemBlock_208 : outputMemBlock_207;
  assign _GEN_1234 = nextBitValid ? outputMemBlock_209 : outputMemBlock_208;
  assign _GEN_1235 = nextBitValid ? outputMemBlock_210 : outputMemBlock_209;
  assign _GEN_1236 = nextBitValid ? outputMemBlock_211 : outputMemBlock_210;
  assign _GEN_1237 = nextBitValid ? outputMemBlock_212 : outputMemBlock_211;
  assign _GEN_1238 = nextBitValid ? outputMemBlock_213 : outputMemBlock_212;
  assign _GEN_1239 = nextBitValid ? outputMemBlock_214 : outputMemBlock_213;
  assign _GEN_1240 = nextBitValid ? outputMemBlock_215 : outputMemBlock_214;
  assign _GEN_1241 = nextBitValid ? outputMemBlock_216 : outputMemBlock_215;
  assign _GEN_1242 = nextBitValid ? outputMemBlock_217 : outputMemBlock_216;
  assign _GEN_1243 = nextBitValid ? outputMemBlock_218 : outputMemBlock_217;
  assign _GEN_1244 = nextBitValid ? outputMemBlock_219 : outputMemBlock_218;
  assign _GEN_1245 = nextBitValid ? outputMemBlock_220 : outputMemBlock_219;
  assign _GEN_1246 = nextBitValid ? outputMemBlock_221 : outputMemBlock_220;
  assign _GEN_1247 = nextBitValid ? outputMemBlock_222 : outputMemBlock_221;
  assign _GEN_1248 = nextBitValid ? outputMemBlock_223 : outputMemBlock_222;
  assign _GEN_1249 = nextBitValid ? outputMemBlock_224 : outputMemBlock_223;
  assign _GEN_1250 = nextBitValid ? outputMemBlock_225 : outputMemBlock_224;
  assign _GEN_1251 = nextBitValid ? outputMemBlock_226 : outputMemBlock_225;
  assign _GEN_1252 = nextBitValid ? outputMemBlock_227 : outputMemBlock_226;
  assign _GEN_1253 = nextBitValid ? outputMemBlock_228 : outputMemBlock_227;
  assign _GEN_1254 = nextBitValid ? outputMemBlock_229 : outputMemBlock_228;
  assign _GEN_1255 = nextBitValid ? outputMemBlock_230 : outputMemBlock_229;
  assign _GEN_1256 = nextBitValid ? outputMemBlock_231 : outputMemBlock_230;
  assign _GEN_1257 = nextBitValid ? outputMemBlock_232 : outputMemBlock_231;
  assign _GEN_1258 = nextBitValid ? outputMemBlock_233 : outputMemBlock_232;
  assign _GEN_1259 = nextBitValid ? outputMemBlock_234 : outputMemBlock_233;
  assign _GEN_1260 = nextBitValid ? outputMemBlock_235 : outputMemBlock_234;
  assign _GEN_1261 = nextBitValid ? outputMemBlock_236 : outputMemBlock_235;
  assign _GEN_1262 = nextBitValid ? outputMemBlock_237 : outputMemBlock_236;
  assign _GEN_1263 = nextBitValid ? outputMemBlock_238 : outputMemBlock_237;
  assign _GEN_1264 = nextBitValid ? outputMemBlock_239 : outputMemBlock_238;
  assign _GEN_1265 = nextBitValid ? outputMemBlock_240 : outputMemBlock_239;
  assign _GEN_1266 = nextBitValid ? outputMemBlock_241 : outputMemBlock_240;
  assign _GEN_1267 = nextBitValid ? outputMemBlock_242 : outputMemBlock_241;
  assign _GEN_1268 = nextBitValid ? outputMemBlock_243 : outputMemBlock_242;
  assign _GEN_1269 = nextBitValid ? outputMemBlock_244 : outputMemBlock_243;
  assign _GEN_1270 = nextBitValid ? outputMemBlock_245 : outputMemBlock_244;
  assign _GEN_1271 = nextBitValid ? outputMemBlock_246 : outputMemBlock_245;
  assign _GEN_1272 = nextBitValid ? outputMemBlock_247 : outputMemBlock_246;
  assign _GEN_1273 = nextBitValid ? outputMemBlock_248 : outputMemBlock_247;
  assign _GEN_1274 = nextBitValid ? outputMemBlock_249 : outputMemBlock_248;
  assign _GEN_1275 = nextBitValid ? outputMemBlock_250 : outputMemBlock_249;
  assign _GEN_1276 = nextBitValid ? outputMemBlock_251 : outputMemBlock_250;
  assign _GEN_1277 = nextBitValid ? outputMemBlock_252 : outputMemBlock_251;
  assign _GEN_1278 = nextBitValid ? outputMemBlock_253 : outputMemBlock_252;
  assign _GEN_1279 = nextBitValid ? outputMemBlock_254 : outputMemBlock_253;
  assign _GEN_1280 = nextBitValid ? outputMemBlock_255 : outputMemBlock_254;
  assign _GEN_1281 = nextBitValid ? outputMemBlock_256 : outputMemBlock_255;
  assign _GEN_1282 = nextBitValid ? outputMemBlock_257 : outputMemBlock_256;
  assign _GEN_1283 = nextBitValid ? outputMemBlock_258 : outputMemBlock_257;
  assign _GEN_1284 = nextBitValid ? outputMemBlock_259 : outputMemBlock_258;
  assign _GEN_1285 = nextBitValid ? outputMemBlock_260 : outputMemBlock_259;
  assign _GEN_1286 = nextBitValid ? outputMemBlock_261 : outputMemBlock_260;
  assign _GEN_1287 = nextBitValid ? outputMemBlock_262 : outputMemBlock_261;
  assign _GEN_1288 = nextBitValid ? outputMemBlock_263 : outputMemBlock_262;
  assign _GEN_1289 = nextBitValid ? outputMemBlock_264 : outputMemBlock_263;
  assign _GEN_1290 = nextBitValid ? outputMemBlock_265 : outputMemBlock_264;
  assign _GEN_1291 = nextBitValid ? outputMemBlock_266 : outputMemBlock_265;
  assign _GEN_1292 = nextBitValid ? outputMemBlock_267 : outputMemBlock_266;
  assign _GEN_1293 = nextBitValid ? outputMemBlock_268 : outputMemBlock_267;
  assign _GEN_1294 = nextBitValid ? outputMemBlock_269 : outputMemBlock_268;
  assign _GEN_1295 = nextBitValid ? outputMemBlock_270 : outputMemBlock_269;
  assign _GEN_1296 = nextBitValid ? outputMemBlock_271 : outputMemBlock_270;
  assign _GEN_1297 = nextBitValid ? outputMemBlock_272 : outputMemBlock_271;
  assign _GEN_1298 = nextBitValid ? outputMemBlock_273 : outputMemBlock_272;
  assign _GEN_1299 = nextBitValid ? outputMemBlock_274 : outputMemBlock_273;
  assign _GEN_1300 = nextBitValid ? outputMemBlock_275 : outputMemBlock_274;
  assign _GEN_1301 = nextBitValid ? outputMemBlock_276 : outputMemBlock_275;
  assign _GEN_1302 = nextBitValid ? outputMemBlock_277 : outputMemBlock_276;
  assign _GEN_1303 = nextBitValid ? outputMemBlock_278 : outputMemBlock_277;
  assign _GEN_1304 = nextBitValid ? outputMemBlock_279 : outputMemBlock_278;
  assign _GEN_1305 = nextBitValid ? outputMemBlock_280 : outputMemBlock_279;
  assign _GEN_1306 = nextBitValid ? outputMemBlock_281 : outputMemBlock_280;
  assign _GEN_1307 = nextBitValid ? outputMemBlock_282 : outputMemBlock_281;
  assign _GEN_1308 = nextBitValid ? outputMemBlock_283 : outputMemBlock_282;
  assign _GEN_1309 = nextBitValid ? outputMemBlock_284 : outputMemBlock_283;
  assign _GEN_1310 = nextBitValid ? outputMemBlock_285 : outputMemBlock_284;
  assign _GEN_1311 = nextBitValid ? outputMemBlock_286 : outputMemBlock_285;
  assign _GEN_1312 = nextBitValid ? outputMemBlock_287 : outputMemBlock_286;
  assign _GEN_1313 = nextBitValid ? outputMemBlock_288 : outputMemBlock_287;
  assign _GEN_1314 = nextBitValid ? outputMemBlock_289 : outputMemBlock_288;
  assign _GEN_1315 = nextBitValid ? outputMemBlock_290 : outputMemBlock_289;
  assign _GEN_1316 = nextBitValid ? outputMemBlock_291 : outputMemBlock_290;
  assign _GEN_1317 = nextBitValid ? outputMemBlock_292 : outputMemBlock_291;
  assign _GEN_1318 = nextBitValid ? outputMemBlock_293 : outputMemBlock_292;
  assign _GEN_1319 = nextBitValid ? outputMemBlock_294 : outputMemBlock_293;
  assign _GEN_1320 = nextBitValid ? outputMemBlock_295 : outputMemBlock_294;
  assign _GEN_1321 = nextBitValid ? outputMemBlock_296 : outputMemBlock_295;
  assign _GEN_1322 = nextBitValid ? outputMemBlock_297 : outputMemBlock_296;
  assign _GEN_1323 = nextBitValid ? outputMemBlock_298 : outputMemBlock_297;
  assign _GEN_1324 = nextBitValid ? outputMemBlock_299 : outputMemBlock_298;
  assign _GEN_1325 = nextBitValid ? outputMemBlock_300 : outputMemBlock_299;
  assign _GEN_1326 = nextBitValid ? outputMemBlock_301 : outputMemBlock_300;
  assign _GEN_1327 = nextBitValid ? outputMemBlock_302 : outputMemBlock_301;
  assign _GEN_1328 = nextBitValid ? outputMemBlock_303 : outputMemBlock_302;
  assign _GEN_1329 = nextBitValid ? outputMemBlock_304 : outputMemBlock_303;
  assign _GEN_1330 = nextBitValid ? outputMemBlock_305 : outputMemBlock_304;
  assign _GEN_1331 = nextBitValid ? outputMemBlock_306 : outputMemBlock_305;
  assign _GEN_1332 = nextBitValid ? outputMemBlock_307 : outputMemBlock_306;
  assign _GEN_1333 = nextBitValid ? outputMemBlock_308 : outputMemBlock_307;
  assign _GEN_1334 = nextBitValid ? outputMemBlock_309 : outputMemBlock_308;
  assign _GEN_1335 = nextBitValid ? outputMemBlock_310 : outputMemBlock_309;
  assign _GEN_1336 = nextBitValid ? outputMemBlock_311 : outputMemBlock_310;
  assign _GEN_1337 = nextBitValid ? outputMemBlock_312 : outputMemBlock_311;
  assign _GEN_1338 = nextBitValid ? outputMemBlock_313 : outputMemBlock_312;
  assign _GEN_1339 = nextBitValid ? outputMemBlock_314 : outputMemBlock_313;
  assign _GEN_1340 = nextBitValid ? outputMemBlock_315 : outputMemBlock_314;
  assign _GEN_1341 = nextBitValid ? outputMemBlock_316 : outputMemBlock_315;
  assign _GEN_1342 = nextBitValid ? outputMemBlock_317 : outputMemBlock_316;
  assign _GEN_1343 = nextBitValid ? outputMemBlock_318 : outputMemBlock_317;
  assign _GEN_1344 = nextBitValid ? outputMemBlock_319 : outputMemBlock_318;
  assign _GEN_1345 = nextBitValid ? outputMemBlock_320 : outputMemBlock_319;
  assign _GEN_1346 = nextBitValid ? outputMemBlock_321 : outputMemBlock_320;
  assign _GEN_1347 = nextBitValid ? outputMemBlock_322 : outputMemBlock_321;
  assign _GEN_1348 = nextBitValid ? outputMemBlock_323 : outputMemBlock_322;
  assign _GEN_1349 = nextBitValid ? outputMemBlock_324 : outputMemBlock_323;
  assign _GEN_1350 = nextBitValid ? outputMemBlock_325 : outputMemBlock_324;
  assign _GEN_1351 = nextBitValid ? outputMemBlock_326 : outputMemBlock_325;
  assign _GEN_1352 = nextBitValid ? outputMemBlock_327 : outputMemBlock_326;
  assign _GEN_1353 = nextBitValid ? outputMemBlock_328 : outputMemBlock_327;
  assign _GEN_1354 = nextBitValid ? outputMemBlock_329 : outputMemBlock_328;
  assign _GEN_1355 = nextBitValid ? outputMemBlock_330 : outputMemBlock_329;
  assign _GEN_1356 = nextBitValid ? outputMemBlock_331 : outputMemBlock_330;
  assign _GEN_1357 = nextBitValid ? outputMemBlock_332 : outputMemBlock_331;
  assign _GEN_1358 = nextBitValid ? outputMemBlock_333 : outputMemBlock_332;
  assign _GEN_1359 = nextBitValid ? outputMemBlock_334 : outputMemBlock_333;
  assign _GEN_1360 = nextBitValid ? outputMemBlock_335 : outputMemBlock_334;
  assign _GEN_1361 = nextBitValid ? outputMemBlock_336 : outputMemBlock_335;
  assign _GEN_1362 = nextBitValid ? outputMemBlock_337 : outputMemBlock_336;
  assign _GEN_1363 = nextBitValid ? outputMemBlock_338 : outputMemBlock_337;
  assign _GEN_1364 = nextBitValid ? outputMemBlock_339 : outputMemBlock_338;
  assign _GEN_1365 = nextBitValid ? outputMemBlock_340 : outputMemBlock_339;
  assign _GEN_1366 = nextBitValid ? outputMemBlock_341 : outputMemBlock_340;
  assign _GEN_1367 = nextBitValid ? outputMemBlock_342 : outputMemBlock_341;
  assign _GEN_1368 = nextBitValid ? outputMemBlock_343 : outputMemBlock_342;
  assign _GEN_1369 = nextBitValid ? outputMemBlock_344 : outputMemBlock_343;
  assign _GEN_1370 = nextBitValid ? outputMemBlock_345 : outputMemBlock_344;
  assign _GEN_1371 = nextBitValid ? outputMemBlock_346 : outputMemBlock_345;
  assign _GEN_1372 = nextBitValid ? outputMemBlock_347 : outputMemBlock_346;
  assign _GEN_1373 = nextBitValid ? outputMemBlock_348 : outputMemBlock_347;
  assign _GEN_1374 = nextBitValid ? outputMemBlock_349 : outputMemBlock_348;
  assign _GEN_1375 = nextBitValid ? outputMemBlock_350 : outputMemBlock_349;
  assign _GEN_1376 = nextBitValid ? outputMemBlock_351 : outputMemBlock_350;
  assign _GEN_1377 = nextBitValid ? outputMemBlock_352 : outputMemBlock_351;
  assign _GEN_1378 = nextBitValid ? outputMemBlock_353 : outputMemBlock_352;
  assign _GEN_1379 = nextBitValid ? outputMemBlock_354 : outputMemBlock_353;
  assign _GEN_1380 = nextBitValid ? outputMemBlock_355 : outputMemBlock_354;
  assign _GEN_1381 = nextBitValid ? outputMemBlock_356 : outputMemBlock_355;
  assign _GEN_1382 = nextBitValid ? outputMemBlock_357 : outputMemBlock_356;
  assign _GEN_1383 = nextBitValid ? outputMemBlock_358 : outputMemBlock_357;
  assign _GEN_1384 = nextBitValid ? outputMemBlock_359 : outputMemBlock_358;
  assign _GEN_1385 = nextBitValid ? outputMemBlock_360 : outputMemBlock_359;
  assign _GEN_1386 = nextBitValid ? outputMemBlock_361 : outputMemBlock_360;
  assign _GEN_1387 = nextBitValid ? outputMemBlock_362 : outputMemBlock_361;
  assign _GEN_1388 = nextBitValid ? outputMemBlock_363 : outputMemBlock_362;
  assign _GEN_1389 = nextBitValid ? outputMemBlock_364 : outputMemBlock_363;
  assign _GEN_1390 = nextBitValid ? outputMemBlock_365 : outputMemBlock_364;
  assign _GEN_1391 = nextBitValid ? outputMemBlock_366 : outputMemBlock_365;
  assign _GEN_1392 = nextBitValid ? outputMemBlock_367 : outputMemBlock_366;
  assign _GEN_1393 = nextBitValid ? outputMemBlock_368 : outputMemBlock_367;
  assign _GEN_1394 = nextBitValid ? outputMemBlock_369 : outputMemBlock_368;
  assign _GEN_1395 = nextBitValid ? outputMemBlock_370 : outputMemBlock_369;
  assign _GEN_1396 = nextBitValid ? outputMemBlock_371 : outputMemBlock_370;
  assign _GEN_1397 = nextBitValid ? outputMemBlock_372 : outputMemBlock_371;
  assign _GEN_1398 = nextBitValid ? outputMemBlock_373 : outputMemBlock_372;
  assign _GEN_1399 = nextBitValid ? outputMemBlock_374 : outputMemBlock_373;
  assign _GEN_1400 = nextBitValid ? outputMemBlock_375 : outputMemBlock_374;
  assign _GEN_1401 = nextBitValid ? outputMemBlock_376 : outputMemBlock_375;
  assign _GEN_1402 = nextBitValid ? outputMemBlock_377 : outputMemBlock_376;
  assign _GEN_1403 = nextBitValid ? outputMemBlock_378 : outputMemBlock_377;
  assign _GEN_1404 = nextBitValid ? outputMemBlock_379 : outputMemBlock_378;
  assign _GEN_1405 = nextBitValid ? outputMemBlock_380 : outputMemBlock_379;
  assign _GEN_1406 = nextBitValid ? outputMemBlock_381 : outputMemBlock_380;
  assign _GEN_1407 = nextBitValid ? outputMemBlock_382 : outputMemBlock_381;
  assign _GEN_1408 = nextBitValid ? outputMemBlock_383 : outputMemBlock_382;
  assign _GEN_1409 = nextBitValid ? outputMemBlock_384 : outputMemBlock_383;
  assign _GEN_1410 = nextBitValid ? outputMemBlock_385 : outputMemBlock_384;
  assign _GEN_1411 = nextBitValid ? outputMemBlock_386 : outputMemBlock_385;
  assign _GEN_1412 = nextBitValid ? outputMemBlock_387 : outputMemBlock_386;
  assign _GEN_1413 = nextBitValid ? outputMemBlock_388 : outputMemBlock_387;
  assign _GEN_1414 = nextBitValid ? outputMemBlock_389 : outputMemBlock_388;
  assign _GEN_1415 = nextBitValid ? outputMemBlock_390 : outputMemBlock_389;
  assign _GEN_1416 = nextBitValid ? outputMemBlock_391 : outputMemBlock_390;
  assign _GEN_1417 = nextBitValid ? outputMemBlock_392 : outputMemBlock_391;
  assign _GEN_1418 = nextBitValid ? outputMemBlock_393 : outputMemBlock_392;
  assign _GEN_1419 = nextBitValid ? outputMemBlock_394 : outputMemBlock_393;
  assign _GEN_1420 = nextBitValid ? outputMemBlock_395 : outputMemBlock_394;
  assign _GEN_1421 = nextBitValid ? outputMemBlock_396 : outputMemBlock_395;
  assign _GEN_1422 = nextBitValid ? outputMemBlock_397 : outputMemBlock_396;
  assign _GEN_1423 = nextBitValid ? outputMemBlock_398 : outputMemBlock_397;
  assign _GEN_1424 = nextBitValid ? outputMemBlock_399 : outputMemBlock_398;
  assign _GEN_1425 = nextBitValid ? outputMemBlock_400 : outputMemBlock_399;
  assign _GEN_1426 = nextBitValid ? outputMemBlock_401 : outputMemBlock_400;
  assign _GEN_1427 = nextBitValid ? outputMemBlock_402 : outputMemBlock_401;
  assign _GEN_1428 = nextBitValid ? outputMemBlock_403 : outputMemBlock_402;
  assign _GEN_1429 = nextBitValid ? outputMemBlock_404 : outputMemBlock_403;
  assign _GEN_1430 = nextBitValid ? outputMemBlock_405 : outputMemBlock_404;
  assign _GEN_1431 = nextBitValid ? outputMemBlock_406 : outputMemBlock_405;
  assign _GEN_1432 = nextBitValid ? outputMemBlock_407 : outputMemBlock_406;
  assign _GEN_1433 = nextBitValid ? outputMemBlock_408 : outputMemBlock_407;
  assign _GEN_1434 = nextBitValid ? outputMemBlock_409 : outputMemBlock_408;
  assign _GEN_1435 = nextBitValid ? outputMemBlock_410 : outputMemBlock_409;
  assign _GEN_1436 = nextBitValid ? outputMemBlock_411 : outputMemBlock_410;
  assign _GEN_1437 = nextBitValid ? outputMemBlock_412 : outputMemBlock_411;
  assign _GEN_1438 = nextBitValid ? outputMemBlock_413 : outputMemBlock_412;
  assign _GEN_1439 = nextBitValid ? outputMemBlock_414 : outputMemBlock_413;
  assign _GEN_1440 = nextBitValid ? outputMemBlock_415 : outputMemBlock_414;
  assign _GEN_1441 = nextBitValid ? outputMemBlock_416 : outputMemBlock_415;
  assign _GEN_1442 = nextBitValid ? outputMemBlock_417 : outputMemBlock_416;
  assign _GEN_1443 = nextBitValid ? outputMemBlock_418 : outputMemBlock_417;
  assign _GEN_1444 = nextBitValid ? outputMemBlock_419 : outputMemBlock_418;
  assign _GEN_1445 = nextBitValid ? outputMemBlock_420 : outputMemBlock_419;
  assign _GEN_1446 = nextBitValid ? outputMemBlock_421 : outputMemBlock_420;
  assign _GEN_1447 = nextBitValid ? outputMemBlock_422 : outputMemBlock_421;
  assign _GEN_1448 = nextBitValid ? outputMemBlock_423 : outputMemBlock_422;
  assign _GEN_1449 = nextBitValid ? outputMemBlock_424 : outputMemBlock_423;
  assign _GEN_1450 = nextBitValid ? outputMemBlock_425 : outputMemBlock_424;
  assign _GEN_1451 = nextBitValid ? outputMemBlock_426 : outputMemBlock_425;
  assign _GEN_1452 = nextBitValid ? outputMemBlock_427 : outputMemBlock_426;
  assign _GEN_1453 = nextBitValid ? outputMemBlock_428 : outputMemBlock_427;
  assign _GEN_1454 = nextBitValid ? outputMemBlock_429 : outputMemBlock_428;
  assign _GEN_1455 = nextBitValid ? outputMemBlock_430 : outputMemBlock_429;
  assign _GEN_1456 = nextBitValid ? outputMemBlock_431 : outputMemBlock_430;
  assign _GEN_1457 = nextBitValid ? outputMemBlock_432 : outputMemBlock_431;
  assign _GEN_1458 = nextBitValid ? outputMemBlock_433 : outputMemBlock_432;
  assign _GEN_1459 = nextBitValid ? outputMemBlock_434 : outputMemBlock_433;
  assign _GEN_1460 = nextBitValid ? outputMemBlock_435 : outputMemBlock_434;
  assign _GEN_1461 = nextBitValid ? outputMemBlock_436 : outputMemBlock_435;
  assign _GEN_1462 = nextBitValid ? outputMemBlock_437 : outputMemBlock_436;
  assign _GEN_1463 = nextBitValid ? outputMemBlock_438 : outputMemBlock_437;
  assign _GEN_1464 = nextBitValid ? outputMemBlock_439 : outputMemBlock_438;
  assign _GEN_1465 = nextBitValid ? outputMemBlock_440 : outputMemBlock_439;
  assign _GEN_1466 = nextBitValid ? outputMemBlock_441 : outputMemBlock_440;
  assign _GEN_1467 = nextBitValid ? outputMemBlock_442 : outputMemBlock_441;
  assign _GEN_1468 = nextBitValid ? outputMemBlock_443 : outputMemBlock_442;
  assign _GEN_1469 = nextBitValid ? outputMemBlock_444 : outputMemBlock_443;
  assign _GEN_1470 = nextBitValid ? outputMemBlock_445 : outputMemBlock_444;
  assign _GEN_1471 = nextBitValid ? outputMemBlock_446 : outputMemBlock_445;
  assign _GEN_1472 = nextBitValid ? outputMemBlock_447 : outputMemBlock_446;
  assign _GEN_1473 = nextBitValid ? outputMemBlock_448 : outputMemBlock_447;
  assign _GEN_1474 = nextBitValid ? outputMemBlock_449 : outputMemBlock_448;
  assign _GEN_1475 = nextBitValid ? outputMemBlock_450 : outputMemBlock_449;
  assign _GEN_1476 = nextBitValid ? outputMemBlock_451 : outputMemBlock_450;
  assign _GEN_1477 = nextBitValid ? outputMemBlock_452 : outputMemBlock_451;
  assign _GEN_1478 = nextBitValid ? outputMemBlock_453 : outputMemBlock_452;
  assign _GEN_1479 = nextBitValid ? outputMemBlock_454 : outputMemBlock_453;
  assign _GEN_1480 = nextBitValid ? outputMemBlock_455 : outputMemBlock_454;
  assign _GEN_1481 = nextBitValid ? outputMemBlock_456 : outputMemBlock_455;
  assign _GEN_1482 = nextBitValid ? outputMemBlock_457 : outputMemBlock_456;
  assign _GEN_1483 = nextBitValid ? outputMemBlock_458 : outputMemBlock_457;
  assign _GEN_1484 = nextBitValid ? outputMemBlock_459 : outputMemBlock_458;
  assign _GEN_1485 = nextBitValid ? outputMemBlock_460 : outputMemBlock_459;
  assign _GEN_1486 = nextBitValid ? outputMemBlock_461 : outputMemBlock_460;
  assign _GEN_1487 = nextBitValid ? outputMemBlock_462 : outputMemBlock_461;
  assign _GEN_1488 = nextBitValid ? outputMemBlock_463 : outputMemBlock_462;
  assign _GEN_1489 = nextBitValid ? outputMemBlock_464 : outputMemBlock_463;
  assign _GEN_1490 = nextBitValid ? outputMemBlock_465 : outputMemBlock_464;
  assign _GEN_1491 = nextBitValid ? outputMemBlock_466 : outputMemBlock_465;
  assign _GEN_1492 = nextBitValid ? outputMemBlock_467 : outputMemBlock_466;
  assign _GEN_1493 = nextBitValid ? outputMemBlock_468 : outputMemBlock_467;
  assign _GEN_1494 = nextBitValid ? outputMemBlock_469 : outputMemBlock_468;
  assign _GEN_1495 = nextBitValid ? outputMemBlock_470 : outputMemBlock_469;
  assign _GEN_1496 = nextBitValid ? outputMemBlock_471 : outputMemBlock_470;
  assign _GEN_1497 = nextBitValid ? outputMemBlock_472 : outputMemBlock_471;
  assign _GEN_1498 = nextBitValid ? outputMemBlock_473 : outputMemBlock_472;
  assign _GEN_1499 = nextBitValid ? outputMemBlock_474 : outputMemBlock_473;
  assign _GEN_1500 = nextBitValid ? outputMemBlock_475 : outputMemBlock_474;
  assign _GEN_1501 = nextBitValid ? outputMemBlock_476 : outputMemBlock_475;
  assign _GEN_1502 = nextBitValid ? outputMemBlock_477 : outputMemBlock_476;
  assign _GEN_1503 = nextBitValid ? outputMemBlock_478 : outputMemBlock_477;
  assign _GEN_1504 = nextBitValid ? outputMemBlock_479 : outputMemBlock_478;
  assign _GEN_1505 = nextBitValid ? outputMemBlock_480 : outputMemBlock_479;
  assign _GEN_1506 = nextBitValid ? outputMemBlock_481 : outputMemBlock_480;
  assign _GEN_1507 = nextBitValid ? outputMemBlock_482 : outputMemBlock_481;
  assign _GEN_1508 = nextBitValid ? outputMemBlock_483 : outputMemBlock_482;
  assign _GEN_1509 = nextBitValid ? outputMemBlock_484 : outputMemBlock_483;
  assign _GEN_1510 = nextBitValid ? outputMemBlock_485 : outputMemBlock_484;
  assign _GEN_1511 = nextBitValid ? outputMemBlock_486 : outputMemBlock_485;
  assign _GEN_1512 = nextBitValid ? outputMemBlock_487 : outputMemBlock_486;
  assign _GEN_1513 = nextBitValid ? outputMemBlock_488 : outputMemBlock_487;
  assign _GEN_1514 = nextBitValid ? outputMemBlock_489 : outputMemBlock_488;
  assign _GEN_1515 = nextBitValid ? outputMemBlock_490 : outputMemBlock_489;
  assign _GEN_1516 = nextBitValid ? outputMemBlock_491 : outputMemBlock_490;
  assign _GEN_1517 = nextBitValid ? outputMemBlock_492 : outputMemBlock_491;
  assign _GEN_1518 = nextBitValid ? outputMemBlock_493 : outputMemBlock_492;
  assign _GEN_1519 = nextBitValid ? outputMemBlock_494 : outputMemBlock_493;
  assign _GEN_1520 = nextBitValid ? outputMemBlock_495 : outputMemBlock_494;
  assign _GEN_1521 = nextBitValid ? outputMemBlock_496 : outputMemBlock_495;
  assign _GEN_1522 = nextBitValid ? outputMemBlock_497 : outputMemBlock_496;
  assign _GEN_1523 = nextBitValid ? outputMemBlock_498 : outputMemBlock_497;
  assign _GEN_1524 = nextBitValid ? outputMemBlock_499 : outputMemBlock_498;
  assign _GEN_1525 = nextBitValid ? outputMemBlock_500 : outputMemBlock_499;
  assign _GEN_1526 = nextBitValid ? outputMemBlock_501 : outputMemBlock_500;
  assign _GEN_1527 = nextBitValid ? outputMemBlock_502 : outputMemBlock_501;
  assign _GEN_1528 = nextBitValid ? outputMemBlock_503 : outputMemBlock_502;
  assign _GEN_1529 = nextBitValid ? outputMemBlock_504 : outputMemBlock_503;
  assign _GEN_1530 = nextBitValid ? outputMemBlock_505 : outputMemBlock_504;
  assign _GEN_1531 = nextBitValid ? outputMemBlock_506 : outputMemBlock_505;
  assign _GEN_1532 = nextBitValid ? outputMemBlock_507 : outputMemBlock_506;
  assign _GEN_1533 = nextBitValid ? outputMemBlock_508 : outputMemBlock_507;
  assign _GEN_1534 = nextBitValid ? outputMemBlock_509 : outputMemBlock_508;
  assign _GEN_1535 = nextBitValid ? outputMemBlock_510 : outputMemBlock_509;
  assign _GEN_1536 = nextBitValid ? outputMemBlock_511 : outputMemBlock_510;
  assign _GEN_1537 = nextBitValid ? _T_1588 : outputBits;
  assign _T_1590 = outputBits == 10'h200;
  assign _T_1593 = io_inputFinished & _T_1053;
  assign _T_1595 = outputBits > 10'h0;
  assign _T_1596 = _T_1593 & _T_1595;
  assign _T_1597 = _T_1590 | _T_1596;
  assign _T_1598 = {outputMemBlock_1,outputMemBlock_0};
  assign _T_1599 = {outputMemBlock_3,outputMemBlock_2};
  assign _T_1600 = {_T_1599,_T_1598};
  assign _T_1601 = {outputMemBlock_5,outputMemBlock_4};
  assign _T_1602 = {outputMemBlock_7,outputMemBlock_6};
  assign _T_1603 = {_T_1602,_T_1601};
  assign _T_1604 = {_T_1603,_T_1600};
  assign _T_1605 = {outputMemBlock_9,outputMemBlock_8};
  assign _T_1606 = {outputMemBlock_11,outputMemBlock_10};
  assign _T_1607 = {_T_1606,_T_1605};
  assign _T_1608 = {outputMemBlock_13,outputMemBlock_12};
  assign _T_1609 = {outputMemBlock_15,outputMemBlock_14};
  assign _T_1610 = {_T_1609,_T_1608};
  assign _T_1611 = {_T_1610,_T_1607};
  assign _T_1612 = {_T_1611,_T_1604};
  assign _T_1613 = {outputMemBlock_17,outputMemBlock_16};
  assign _T_1614 = {outputMemBlock_19,outputMemBlock_18};
  assign _T_1615 = {_T_1614,_T_1613};
  assign _T_1616 = {outputMemBlock_21,outputMemBlock_20};
  assign _T_1617 = {outputMemBlock_23,outputMemBlock_22};
  assign _T_1618 = {_T_1617,_T_1616};
  assign _T_1619 = {_T_1618,_T_1615};
  assign _T_1620 = {outputMemBlock_25,outputMemBlock_24};
  assign _T_1621 = {outputMemBlock_27,outputMemBlock_26};
  assign _T_1622 = {_T_1621,_T_1620};
  assign _T_1623 = {outputMemBlock_29,outputMemBlock_28};
  assign _T_1624 = {outputMemBlock_31,outputMemBlock_30};
  assign _T_1625 = {_T_1624,_T_1623};
  assign _T_1626 = {_T_1625,_T_1622};
  assign _T_1627 = {_T_1626,_T_1619};
  assign _T_1628 = {_T_1627,_T_1612};
  assign _T_1629 = {outputMemBlock_33,outputMemBlock_32};
  assign _T_1630 = {outputMemBlock_35,outputMemBlock_34};
  assign _T_1631 = {_T_1630,_T_1629};
  assign _T_1632 = {outputMemBlock_37,outputMemBlock_36};
  assign _T_1633 = {outputMemBlock_39,outputMemBlock_38};
  assign _T_1634 = {_T_1633,_T_1632};
  assign _T_1635 = {_T_1634,_T_1631};
  assign _T_1636 = {outputMemBlock_41,outputMemBlock_40};
  assign _T_1637 = {outputMemBlock_43,outputMemBlock_42};
  assign _T_1638 = {_T_1637,_T_1636};
  assign _T_1639 = {outputMemBlock_45,outputMemBlock_44};
  assign _T_1640 = {outputMemBlock_47,outputMemBlock_46};
  assign _T_1641 = {_T_1640,_T_1639};
  assign _T_1642 = {_T_1641,_T_1638};
  assign _T_1643 = {_T_1642,_T_1635};
  assign _T_1644 = {outputMemBlock_49,outputMemBlock_48};
  assign _T_1645 = {outputMemBlock_51,outputMemBlock_50};
  assign _T_1646 = {_T_1645,_T_1644};
  assign _T_1647 = {outputMemBlock_53,outputMemBlock_52};
  assign _T_1648 = {outputMemBlock_55,outputMemBlock_54};
  assign _T_1649 = {_T_1648,_T_1647};
  assign _T_1650 = {_T_1649,_T_1646};
  assign _T_1651 = {outputMemBlock_57,outputMemBlock_56};
  assign _T_1652 = {outputMemBlock_59,outputMemBlock_58};
  assign _T_1653 = {_T_1652,_T_1651};
  assign _T_1654 = {outputMemBlock_61,outputMemBlock_60};
  assign _T_1655 = {outputMemBlock_63,outputMemBlock_62};
  assign _T_1656 = {_T_1655,_T_1654};
  assign _T_1657 = {_T_1656,_T_1653};
  assign _T_1658 = {_T_1657,_T_1650};
  assign _T_1659 = {_T_1658,_T_1643};
  assign _T_1660 = {_T_1659,_T_1628};
  assign _T_1661 = {outputMemBlock_65,outputMemBlock_64};
  assign _T_1662 = {outputMemBlock_67,outputMemBlock_66};
  assign _T_1663 = {_T_1662,_T_1661};
  assign _T_1664 = {outputMemBlock_69,outputMemBlock_68};
  assign _T_1665 = {outputMemBlock_71,outputMemBlock_70};
  assign _T_1666 = {_T_1665,_T_1664};
  assign _T_1667 = {_T_1666,_T_1663};
  assign _T_1668 = {outputMemBlock_73,outputMemBlock_72};
  assign _T_1669 = {outputMemBlock_75,outputMemBlock_74};
  assign _T_1670 = {_T_1669,_T_1668};
  assign _T_1671 = {outputMemBlock_77,outputMemBlock_76};
  assign _T_1672 = {outputMemBlock_79,outputMemBlock_78};
  assign _T_1673 = {_T_1672,_T_1671};
  assign _T_1674 = {_T_1673,_T_1670};
  assign _T_1675 = {_T_1674,_T_1667};
  assign _T_1676 = {outputMemBlock_81,outputMemBlock_80};
  assign _T_1677 = {outputMemBlock_83,outputMemBlock_82};
  assign _T_1678 = {_T_1677,_T_1676};
  assign _T_1679 = {outputMemBlock_85,outputMemBlock_84};
  assign _T_1680 = {outputMemBlock_87,outputMemBlock_86};
  assign _T_1681 = {_T_1680,_T_1679};
  assign _T_1682 = {_T_1681,_T_1678};
  assign _T_1683 = {outputMemBlock_89,outputMemBlock_88};
  assign _T_1684 = {outputMemBlock_91,outputMemBlock_90};
  assign _T_1685 = {_T_1684,_T_1683};
  assign _T_1686 = {outputMemBlock_93,outputMemBlock_92};
  assign _T_1687 = {outputMemBlock_95,outputMemBlock_94};
  assign _T_1688 = {_T_1687,_T_1686};
  assign _T_1689 = {_T_1688,_T_1685};
  assign _T_1690 = {_T_1689,_T_1682};
  assign _T_1691 = {_T_1690,_T_1675};
  assign _T_1692 = {outputMemBlock_97,outputMemBlock_96};
  assign _T_1693 = {outputMemBlock_99,outputMemBlock_98};
  assign _T_1694 = {_T_1693,_T_1692};
  assign _T_1695 = {outputMemBlock_101,outputMemBlock_100};
  assign _T_1696 = {outputMemBlock_103,outputMemBlock_102};
  assign _T_1697 = {_T_1696,_T_1695};
  assign _T_1698 = {_T_1697,_T_1694};
  assign _T_1699 = {outputMemBlock_105,outputMemBlock_104};
  assign _T_1700 = {outputMemBlock_107,outputMemBlock_106};
  assign _T_1701 = {_T_1700,_T_1699};
  assign _T_1702 = {outputMemBlock_109,outputMemBlock_108};
  assign _T_1703 = {outputMemBlock_111,outputMemBlock_110};
  assign _T_1704 = {_T_1703,_T_1702};
  assign _T_1705 = {_T_1704,_T_1701};
  assign _T_1706 = {_T_1705,_T_1698};
  assign _T_1707 = {outputMemBlock_113,outputMemBlock_112};
  assign _T_1708 = {outputMemBlock_115,outputMemBlock_114};
  assign _T_1709 = {_T_1708,_T_1707};
  assign _T_1710 = {outputMemBlock_117,outputMemBlock_116};
  assign _T_1711 = {outputMemBlock_119,outputMemBlock_118};
  assign _T_1712 = {_T_1711,_T_1710};
  assign _T_1713 = {_T_1712,_T_1709};
  assign _T_1714 = {outputMemBlock_121,outputMemBlock_120};
  assign _T_1715 = {outputMemBlock_123,outputMemBlock_122};
  assign _T_1716 = {_T_1715,_T_1714};
  assign _T_1717 = {outputMemBlock_125,outputMemBlock_124};
  assign _T_1718 = {outputMemBlock_127,outputMemBlock_126};
  assign _T_1719 = {_T_1718,_T_1717};
  assign _T_1720 = {_T_1719,_T_1716};
  assign _T_1721 = {_T_1720,_T_1713};
  assign _T_1722 = {_T_1721,_T_1706};
  assign _T_1723 = {_T_1722,_T_1691};
  assign _T_1724 = {_T_1723,_T_1660};
  assign _T_1725 = {outputMemBlock_129,outputMemBlock_128};
  assign _T_1726 = {outputMemBlock_131,outputMemBlock_130};
  assign _T_1727 = {_T_1726,_T_1725};
  assign _T_1728 = {outputMemBlock_133,outputMemBlock_132};
  assign _T_1729 = {outputMemBlock_135,outputMemBlock_134};
  assign _T_1730 = {_T_1729,_T_1728};
  assign _T_1731 = {_T_1730,_T_1727};
  assign _T_1732 = {outputMemBlock_137,outputMemBlock_136};
  assign _T_1733 = {outputMemBlock_139,outputMemBlock_138};
  assign _T_1734 = {_T_1733,_T_1732};
  assign _T_1735 = {outputMemBlock_141,outputMemBlock_140};
  assign _T_1736 = {outputMemBlock_143,outputMemBlock_142};
  assign _T_1737 = {_T_1736,_T_1735};
  assign _T_1738 = {_T_1737,_T_1734};
  assign _T_1739 = {_T_1738,_T_1731};
  assign _T_1740 = {outputMemBlock_145,outputMemBlock_144};
  assign _T_1741 = {outputMemBlock_147,outputMemBlock_146};
  assign _T_1742 = {_T_1741,_T_1740};
  assign _T_1743 = {outputMemBlock_149,outputMemBlock_148};
  assign _T_1744 = {outputMemBlock_151,outputMemBlock_150};
  assign _T_1745 = {_T_1744,_T_1743};
  assign _T_1746 = {_T_1745,_T_1742};
  assign _T_1747 = {outputMemBlock_153,outputMemBlock_152};
  assign _T_1748 = {outputMemBlock_155,outputMemBlock_154};
  assign _T_1749 = {_T_1748,_T_1747};
  assign _T_1750 = {outputMemBlock_157,outputMemBlock_156};
  assign _T_1751 = {outputMemBlock_159,outputMemBlock_158};
  assign _T_1752 = {_T_1751,_T_1750};
  assign _T_1753 = {_T_1752,_T_1749};
  assign _T_1754 = {_T_1753,_T_1746};
  assign _T_1755 = {_T_1754,_T_1739};
  assign _T_1756 = {outputMemBlock_161,outputMemBlock_160};
  assign _T_1757 = {outputMemBlock_163,outputMemBlock_162};
  assign _T_1758 = {_T_1757,_T_1756};
  assign _T_1759 = {outputMemBlock_165,outputMemBlock_164};
  assign _T_1760 = {outputMemBlock_167,outputMemBlock_166};
  assign _T_1761 = {_T_1760,_T_1759};
  assign _T_1762 = {_T_1761,_T_1758};
  assign _T_1763 = {outputMemBlock_169,outputMemBlock_168};
  assign _T_1764 = {outputMemBlock_171,outputMemBlock_170};
  assign _T_1765 = {_T_1764,_T_1763};
  assign _T_1766 = {outputMemBlock_173,outputMemBlock_172};
  assign _T_1767 = {outputMemBlock_175,outputMemBlock_174};
  assign _T_1768 = {_T_1767,_T_1766};
  assign _T_1769 = {_T_1768,_T_1765};
  assign _T_1770 = {_T_1769,_T_1762};
  assign _T_1771 = {outputMemBlock_177,outputMemBlock_176};
  assign _T_1772 = {outputMemBlock_179,outputMemBlock_178};
  assign _T_1773 = {_T_1772,_T_1771};
  assign _T_1774 = {outputMemBlock_181,outputMemBlock_180};
  assign _T_1775 = {outputMemBlock_183,outputMemBlock_182};
  assign _T_1776 = {_T_1775,_T_1774};
  assign _T_1777 = {_T_1776,_T_1773};
  assign _T_1778 = {outputMemBlock_185,outputMemBlock_184};
  assign _T_1779 = {outputMemBlock_187,outputMemBlock_186};
  assign _T_1780 = {_T_1779,_T_1778};
  assign _T_1781 = {outputMemBlock_189,outputMemBlock_188};
  assign _T_1782 = {outputMemBlock_191,outputMemBlock_190};
  assign _T_1783 = {_T_1782,_T_1781};
  assign _T_1784 = {_T_1783,_T_1780};
  assign _T_1785 = {_T_1784,_T_1777};
  assign _T_1786 = {_T_1785,_T_1770};
  assign _T_1787 = {_T_1786,_T_1755};
  assign _T_1788 = {outputMemBlock_193,outputMemBlock_192};
  assign _T_1789 = {outputMemBlock_195,outputMemBlock_194};
  assign _T_1790 = {_T_1789,_T_1788};
  assign _T_1791 = {outputMemBlock_197,outputMemBlock_196};
  assign _T_1792 = {outputMemBlock_199,outputMemBlock_198};
  assign _T_1793 = {_T_1792,_T_1791};
  assign _T_1794 = {_T_1793,_T_1790};
  assign _T_1795 = {outputMemBlock_201,outputMemBlock_200};
  assign _T_1796 = {outputMemBlock_203,outputMemBlock_202};
  assign _T_1797 = {_T_1796,_T_1795};
  assign _T_1798 = {outputMemBlock_205,outputMemBlock_204};
  assign _T_1799 = {outputMemBlock_207,outputMemBlock_206};
  assign _T_1800 = {_T_1799,_T_1798};
  assign _T_1801 = {_T_1800,_T_1797};
  assign _T_1802 = {_T_1801,_T_1794};
  assign _T_1803 = {outputMemBlock_209,outputMemBlock_208};
  assign _T_1804 = {outputMemBlock_211,outputMemBlock_210};
  assign _T_1805 = {_T_1804,_T_1803};
  assign _T_1806 = {outputMemBlock_213,outputMemBlock_212};
  assign _T_1807 = {outputMemBlock_215,outputMemBlock_214};
  assign _T_1808 = {_T_1807,_T_1806};
  assign _T_1809 = {_T_1808,_T_1805};
  assign _T_1810 = {outputMemBlock_217,outputMemBlock_216};
  assign _T_1811 = {outputMemBlock_219,outputMemBlock_218};
  assign _T_1812 = {_T_1811,_T_1810};
  assign _T_1813 = {outputMemBlock_221,outputMemBlock_220};
  assign _T_1814 = {outputMemBlock_223,outputMemBlock_222};
  assign _T_1815 = {_T_1814,_T_1813};
  assign _T_1816 = {_T_1815,_T_1812};
  assign _T_1817 = {_T_1816,_T_1809};
  assign _T_1818 = {_T_1817,_T_1802};
  assign _T_1819 = {outputMemBlock_225,outputMemBlock_224};
  assign _T_1820 = {outputMemBlock_227,outputMemBlock_226};
  assign _T_1821 = {_T_1820,_T_1819};
  assign _T_1822 = {outputMemBlock_229,outputMemBlock_228};
  assign _T_1823 = {outputMemBlock_231,outputMemBlock_230};
  assign _T_1824 = {_T_1823,_T_1822};
  assign _T_1825 = {_T_1824,_T_1821};
  assign _T_1826 = {outputMemBlock_233,outputMemBlock_232};
  assign _T_1827 = {outputMemBlock_235,outputMemBlock_234};
  assign _T_1828 = {_T_1827,_T_1826};
  assign _T_1829 = {outputMemBlock_237,outputMemBlock_236};
  assign _T_1830 = {outputMemBlock_239,outputMemBlock_238};
  assign _T_1831 = {_T_1830,_T_1829};
  assign _T_1832 = {_T_1831,_T_1828};
  assign _T_1833 = {_T_1832,_T_1825};
  assign _T_1834 = {outputMemBlock_241,outputMemBlock_240};
  assign _T_1835 = {outputMemBlock_243,outputMemBlock_242};
  assign _T_1836 = {_T_1835,_T_1834};
  assign _T_1837 = {outputMemBlock_245,outputMemBlock_244};
  assign _T_1838 = {outputMemBlock_247,outputMemBlock_246};
  assign _T_1839 = {_T_1838,_T_1837};
  assign _T_1840 = {_T_1839,_T_1836};
  assign _T_1841 = {outputMemBlock_249,outputMemBlock_248};
  assign _T_1842 = {outputMemBlock_251,outputMemBlock_250};
  assign _T_1843 = {_T_1842,_T_1841};
  assign _T_1844 = {outputMemBlock_253,outputMemBlock_252};
  assign _T_1845 = {outputMemBlock_255,outputMemBlock_254};
  assign _T_1846 = {_T_1845,_T_1844};
  assign _T_1847 = {_T_1846,_T_1843};
  assign _T_1848 = {_T_1847,_T_1840};
  assign _T_1849 = {_T_1848,_T_1833};
  assign _T_1850 = {_T_1849,_T_1818};
  assign _T_1851 = {_T_1850,_T_1787};
  assign _T_1852 = {_T_1851,_T_1724};
  assign _T_1853 = {outputMemBlock_257,outputMemBlock_256};
  assign _T_1854 = {outputMemBlock_259,outputMemBlock_258};
  assign _T_1855 = {_T_1854,_T_1853};
  assign _T_1856 = {outputMemBlock_261,outputMemBlock_260};
  assign _T_1857 = {outputMemBlock_263,outputMemBlock_262};
  assign _T_1858 = {_T_1857,_T_1856};
  assign _T_1859 = {_T_1858,_T_1855};
  assign _T_1860 = {outputMemBlock_265,outputMemBlock_264};
  assign _T_1861 = {outputMemBlock_267,outputMemBlock_266};
  assign _T_1862 = {_T_1861,_T_1860};
  assign _T_1863 = {outputMemBlock_269,outputMemBlock_268};
  assign _T_1864 = {outputMemBlock_271,outputMemBlock_270};
  assign _T_1865 = {_T_1864,_T_1863};
  assign _T_1866 = {_T_1865,_T_1862};
  assign _T_1867 = {_T_1866,_T_1859};
  assign _T_1868 = {outputMemBlock_273,outputMemBlock_272};
  assign _T_1869 = {outputMemBlock_275,outputMemBlock_274};
  assign _T_1870 = {_T_1869,_T_1868};
  assign _T_1871 = {outputMemBlock_277,outputMemBlock_276};
  assign _T_1872 = {outputMemBlock_279,outputMemBlock_278};
  assign _T_1873 = {_T_1872,_T_1871};
  assign _T_1874 = {_T_1873,_T_1870};
  assign _T_1875 = {outputMemBlock_281,outputMemBlock_280};
  assign _T_1876 = {outputMemBlock_283,outputMemBlock_282};
  assign _T_1877 = {_T_1876,_T_1875};
  assign _T_1878 = {outputMemBlock_285,outputMemBlock_284};
  assign _T_1879 = {outputMemBlock_287,outputMemBlock_286};
  assign _T_1880 = {_T_1879,_T_1878};
  assign _T_1881 = {_T_1880,_T_1877};
  assign _T_1882 = {_T_1881,_T_1874};
  assign _T_1883 = {_T_1882,_T_1867};
  assign _T_1884 = {outputMemBlock_289,outputMemBlock_288};
  assign _T_1885 = {outputMemBlock_291,outputMemBlock_290};
  assign _T_1886 = {_T_1885,_T_1884};
  assign _T_1887 = {outputMemBlock_293,outputMemBlock_292};
  assign _T_1888 = {outputMemBlock_295,outputMemBlock_294};
  assign _T_1889 = {_T_1888,_T_1887};
  assign _T_1890 = {_T_1889,_T_1886};
  assign _T_1891 = {outputMemBlock_297,outputMemBlock_296};
  assign _T_1892 = {outputMemBlock_299,outputMemBlock_298};
  assign _T_1893 = {_T_1892,_T_1891};
  assign _T_1894 = {outputMemBlock_301,outputMemBlock_300};
  assign _T_1895 = {outputMemBlock_303,outputMemBlock_302};
  assign _T_1896 = {_T_1895,_T_1894};
  assign _T_1897 = {_T_1896,_T_1893};
  assign _T_1898 = {_T_1897,_T_1890};
  assign _T_1899 = {outputMemBlock_305,outputMemBlock_304};
  assign _T_1900 = {outputMemBlock_307,outputMemBlock_306};
  assign _T_1901 = {_T_1900,_T_1899};
  assign _T_1902 = {outputMemBlock_309,outputMemBlock_308};
  assign _T_1903 = {outputMemBlock_311,outputMemBlock_310};
  assign _T_1904 = {_T_1903,_T_1902};
  assign _T_1905 = {_T_1904,_T_1901};
  assign _T_1906 = {outputMemBlock_313,outputMemBlock_312};
  assign _T_1907 = {outputMemBlock_315,outputMemBlock_314};
  assign _T_1908 = {_T_1907,_T_1906};
  assign _T_1909 = {outputMemBlock_317,outputMemBlock_316};
  assign _T_1910 = {outputMemBlock_319,outputMemBlock_318};
  assign _T_1911 = {_T_1910,_T_1909};
  assign _T_1912 = {_T_1911,_T_1908};
  assign _T_1913 = {_T_1912,_T_1905};
  assign _T_1914 = {_T_1913,_T_1898};
  assign _T_1915 = {_T_1914,_T_1883};
  assign _T_1916 = {outputMemBlock_321,outputMemBlock_320};
  assign _T_1917 = {outputMemBlock_323,outputMemBlock_322};
  assign _T_1918 = {_T_1917,_T_1916};
  assign _T_1919 = {outputMemBlock_325,outputMemBlock_324};
  assign _T_1920 = {outputMemBlock_327,outputMemBlock_326};
  assign _T_1921 = {_T_1920,_T_1919};
  assign _T_1922 = {_T_1921,_T_1918};
  assign _T_1923 = {outputMemBlock_329,outputMemBlock_328};
  assign _T_1924 = {outputMemBlock_331,outputMemBlock_330};
  assign _T_1925 = {_T_1924,_T_1923};
  assign _T_1926 = {outputMemBlock_333,outputMemBlock_332};
  assign _T_1927 = {outputMemBlock_335,outputMemBlock_334};
  assign _T_1928 = {_T_1927,_T_1926};
  assign _T_1929 = {_T_1928,_T_1925};
  assign _T_1930 = {_T_1929,_T_1922};
  assign _T_1931 = {outputMemBlock_337,outputMemBlock_336};
  assign _T_1932 = {outputMemBlock_339,outputMemBlock_338};
  assign _T_1933 = {_T_1932,_T_1931};
  assign _T_1934 = {outputMemBlock_341,outputMemBlock_340};
  assign _T_1935 = {outputMemBlock_343,outputMemBlock_342};
  assign _T_1936 = {_T_1935,_T_1934};
  assign _T_1937 = {_T_1936,_T_1933};
  assign _T_1938 = {outputMemBlock_345,outputMemBlock_344};
  assign _T_1939 = {outputMemBlock_347,outputMemBlock_346};
  assign _T_1940 = {_T_1939,_T_1938};
  assign _T_1941 = {outputMemBlock_349,outputMemBlock_348};
  assign _T_1942 = {outputMemBlock_351,outputMemBlock_350};
  assign _T_1943 = {_T_1942,_T_1941};
  assign _T_1944 = {_T_1943,_T_1940};
  assign _T_1945 = {_T_1944,_T_1937};
  assign _T_1946 = {_T_1945,_T_1930};
  assign _T_1947 = {outputMemBlock_353,outputMemBlock_352};
  assign _T_1948 = {outputMemBlock_355,outputMemBlock_354};
  assign _T_1949 = {_T_1948,_T_1947};
  assign _T_1950 = {outputMemBlock_357,outputMemBlock_356};
  assign _T_1951 = {outputMemBlock_359,outputMemBlock_358};
  assign _T_1952 = {_T_1951,_T_1950};
  assign _T_1953 = {_T_1952,_T_1949};
  assign _T_1954 = {outputMemBlock_361,outputMemBlock_360};
  assign _T_1955 = {outputMemBlock_363,outputMemBlock_362};
  assign _T_1956 = {_T_1955,_T_1954};
  assign _T_1957 = {outputMemBlock_365,outputMemBlock_364};
  assign _T_1958 = {outputMemBlock_367,outputMemBlock_366};
  assign _T_1959 = {_T_1958,_T_1957};
  assign _T_1960 = {_T_1959,_T_1956};
  assign _T_1961 = {_T_1960,_T_1953};
  assign _T_1962 = {outputMemBlock_369,outputMemBlock_368};
  assign _T_1963 = {outputMemBlock_371,outputMemBlock_370};
  assign _T_1964 = {_T_1963,_T_1962};
  assign _T_1965 = {outputMemBlock_373,outputMemBlock_372};
  assign _T_1966 = {outputMemBlock_375,outputMemBlock_374};
  assign _T_1967 = {_T_1966,_T_1965};
  assign _T_1968 = {_T_1967,_T_1964};
  assign _T_1969 = {outputMemBlock_377,outputMemBlock_376};
  assign _T_1970 = {outputMemBlock_379,outputMemBlock_378};
  assign _T_1971 = {_T_1970,_T_1969};
  assign _T_1972 = {outputMemBlock_381,outputMemBlock_380};
  assign _T_1973 = {outputMemBlock_383,outputMemBlock_382};
  assign _T_1974 = {_T_1973,_T_1972};
  assign _T_1975 = {_T_1974,_T_1971};
  assign _T_1976 = {_T_1975,_T_1968};
  assign _T_1977 = {_T_1976,_T_1961};
  assign _T_1978 = {_T_1977,_T_1946};
  assign _T_1979 = {_T_1978,_T_1915};
  assign _T_1980 = {outputMemBlock_385,outputMemBlock_384};
  assign _T_1981 = {outputMemBlock_387,outputMemBlock_386};
  assign _T_1982 = {_T_1981,_T_1980};
  assign _T_1983 = {outputMemBlock_389,outputMemBlock_388};
  assign _T_1984 = {outputMemBlock_391,outputMemBlock_390};
  assign _T_1985 = {_T_1984,_T_1983};
  assign _T_1986 = {_T_1985,_T_1982};
  assign _T_1987 = {outputMemBlock_393,outputMemBlock_392};
  assign _T_1988 = {outputMemBlock_395,outputMemBlock_394};
  assign _T_1989 = {_T_1988,_T_1987};
  assign _T_1990 = {outputMemBlock_397,outputMemBlock_396};
  assign _T_1991 = {outputMemBlock_399,outputMemBlock_398};
  assign _T_1992 = {_T_1991,_T_1990};
  assign _T_1993 = {_T_1992,_T_1989};
  assign _T_1994 = {_T_1993,_T_1986};
  assign _T_1995 = {outputMemBlock_401,outputMemBlock_400};
  assign _T_1996 = {outputMemBlock_403,outputMemBlock_402};
  assign _T_1997 = {_T_1996,_T_1995};
  assign _T_1998 = {outputMemBlock_405,outputMemBlock_404};
  assign _T_1999 = {outputMemBlock_407,outputMemBlock_406};
  assign _T_2000 = {_T_1999,_T_1998};
  assign _T_2001 = {_T_2000,_T_1997};
  assign _T_2002 = {outputMemBlock_409,outputMemBlock_408};
  assign _T_2003 = {outputMemBlock_411,outputMemBlock_410};
  assign _T_2004 = {_T_2003,_T_2002};
  assign _T_2005 = {outputMemBlock_413,outputMemBlock_412};
  assign _T_2006 = {outputMemBlock_415,outputMemBlock_414};
  assign _T_2007 = {_T_2006,_T_2005};
  assign _T_2008 = {_T_2007,_T_2004};
  assign _T_2009 = {_T_2008,_T_2001};
  assign _T_2010 = {_T_2009,_T_1994};
  assign _T_2011 = {outputMemBlock_417,outputMemBlock_416};
  assign _T_2012 = {outputMemBlock_419,outputMemBlock_418};
  assign _T_2013 = {_T_2012,_T_2011};
  assign _T_2014 = {outputMemBlock_421,outputMemBlock_420};
  assign _T_2015 = {outputMemBlock_423,outputMemBlock_422};
  assign _T_2016 = {_T_2015,_T_2014};
  assign _T_2017 = {_T_2016,_T_2013};
  assign _T_2018 = {outputMemBlock_425,outputMemBlock_424};
  assign _T_2019 = {outputMemBlock_427,outputMemBlock_426};
  assign _T_2020 = {_T_2019,_T_2018};
  assign _T_2021 = {outputMemBlock_429,outputMemBlock_428};
  assign _T_2022 = {outputMemBlock_431,outputMemBlock_430};
  assign _T_2023 = {_T_2022,_T_2021};
  assign _T_2024 = {_T_2023,_T_2020};
  assign _T_2025 = {_T_2024,_T_2017};
  assign _T_2026 = {outputMemBlock_433,outputMemBlock_432};
  assign _T_2027 = {outputMemBlock_435,outputMemBlock_434};
  assign _T_2028 = {_T_2027,_T_2026};
  assign _T_2029 = {outputMemBlock_437,outputMemBlock_436};
  assign _T_2030 = {outputMemBlock_439,outputMemBlock_438};
  assign _T_2031 = {_T_2030,_T_2029};
  assign _T_2032 = {_T_2031,_T_2028};
  assign _T_2033 = {outputMemBlock_441,outputMemBlock_440};
  assign _T_2034 = {outputMemBlock_443,outputMemBlock_442};
  assign _T_2035 = {_T_2034,_T_2033};
  assign _T_2036 = {outputMemBlock_445,outputMemBlock_444};
  assign _T_2037 = {outputMemBlock_447,outputMemBlock_446};
  assign _T_2038 = {_T_2037,_T_2036};
  assign _T_2039 = {_T_2038,_T_2035};
  assign _T_2040 = {_T_2039,_T_2032};
  assign _T_2041 = {_T_2040,_T_2025};
  assign _T_2042 = {_T_2041,_T_2010};
  assign _T_2043 = {outputMemBlock_449,outputMemBlock_448};
  assign _T_2044 = {outputMemBlock_451,outputMemBlock_450};
  assign _T_2045 = {_T_2044,_T_2043};
  assign _T_2046 = {outputMemBlock_453,outputMemBlock_452};
  assign _T_2047 = {outputMemBlock_455,outputMemBlock_454};
  assign _T_2048 = {_T_2047,_T_2046};
  assign _T_2049 = {_T_2048,_T_2045};
  assign _T_2050 = {outputMemBlock_457,outputMemBlock_456};
  assign _T_2051 = {outputMemBlock_459,outputMemBlock_458};
  assign _T_2052 = {_T_2051,_T_2050};
  assign _T_2053 = {outputMemBlock_461,outputMemBlock_460};
  assign _T_2054 = {outputMemBlock_463,outputMemBlock_462};
  assign _T_2055 = {_T_2054,_T_2053};
  assign _T_2056 = {_T_2055,_T_2052};
  assign _T_2057 = {_T_2056,_T_2049};
  assign _T_2058 = {outputMemBlock_465,outputMemBlock_464};
  assign _T_2059 = {outputMemBlock_467,outputMemBlock_466};
  assign _T_2060 = {_T_2059,_T_2058};
  assign _T_2061 = {outputMemBlock_469,outputMemBlock_468};
  assign _T_2062 = {outputMemBlock_471,outputMemBlock_470};
  assign _T_2063 = {_T_2062,_T_2061};
  assign _T_2064 = {_T_2063,_T_2060};
  assign _T_2065 = {outputMemBlock_473,outputMemBlock_472};
  assign _T_2066 = {outputMemBlock_475,outputMemBlock_474};
  assign _T_2067 = {_T_2066,_T_2065};
  assign _T_2068 = {outputMemBlock_477,outputMemBlock_476};
  assign _T_2069 = {outputMemBlock_479,outputMemBlock_478};
  assign _T_2070 = {_T_2069,_T_2068};
  assign _T_2071 = {_T_2070,_T_2067};
  assign _T_2072 = {_T_2071,_T_2064};
  assign _T_2073 = {_T_2072,_T_2057};
  assign _T_2074 = {outputMemBlock_481,outputMemBlock_480};
  assign _T_2075 = {outputMemBlock_483,outputMemBlock_482};
  assign _T_2076 = {_T_2075,_T_2074};
  assign _T_2077 = {outputMemBlock_485,outputMemBlock_484};
  assign _T_2078 = {outputMemBlock_487,outputMemBlock_486};
  assign _T_2079 = {_T_2078,_T_2077};
  assign _T_2080 = {_T_2079,_T_2076};
  assign _T_2081 = {outputMemBlock_489,outputMemBlock_488};
  assign _T_2082 = {outputMemBlock_491,outputMemBlock_490};
  assign _T_2083 = {_T_2082,_T_2081};
  assign _T_2084 = {outputMemBlock_493,outputMemBlock_492};
  assign _T_2085 = {outputMemBlock_495,outputMemBlock_494};
  assign _T_2086 = {_T_2085,_T_2084};
  assign _T_2087 = {_T_2086,_T_2083};
  assign _T_2088 = {_T_2087,_T_2080};
  assign _T_2089 = {outputMemBlock_497,outputMemBlock_496};
  assign _T_2090 = {outputMemBlock_499,outputMemBlock_498};
  assign _T_2091 = {_T_2090,_T_2089};
  assign _T_2092 = {outputMemBlock_501,outputMemBlock_500};
  assign _T_2093 = {outputMemBlock_503,outputMemBlock_502};
  assign _T_2094 = {_T_2093,_T_2092};
  assign _T_2095 = {_T_2094,_T_2091};
  assign _T_2096 = {outputMemBlock_505,outputMemBlock_504};
  assign _T_2097 = {outputMemBlock_507,outputMemBlock_506};
  assign _T_2098 = {_T_2097,_T_2096};
  assign _T_2099 = {outputMemBlock_509,outputMemBlock_508};
  assign _T_2100 = {outputMemBlock_511,outputMemBlock_510};
  assign _T_2101 = {_T_2100,_T_2099};
  assign _T_2102 = {_T_2101,_T_2098};
  assign _T_2103 = {_T_2102,_T_2095};
  assign _T_2104 = {_T_2103,_T_2088};
  assign _T_2105 = {_T_2104,_T_2073};
  assign _T_2106 = {_T_2105,_T_2042};
  assign _T_2107 = {_T_2106,_T_1979};
  assign _T_2108 = {_T_2107,_T_1852};
  assign _T_2113 = outputBits == 10'h0;
  assign _T_2114 = _T_1593 & _T_2113;
  assign _GEN_1538 = io_outputMemFlushed ? 10'h0 : _GEN_1537;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1539 = {1{$random}};
  inputMemBlock_0 = _GEN_1539[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1540 = {1{$random}};
  inputMemBlock_1 = _GEN_1540[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1541 = {1{$random}};
  inputMemBlock_2 = _GEN_1541[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1542 = {1{$random}};
  inputMemBlock_3 = _GEN_1542[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1543 = {1{$random}};
  inputMemBlock_4 = _GEN_1543[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1544 = {1{$random}};
  inputMemBlock_5 = _GEN_1544[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1545 = {1{$random}};
  inputMemBlock_6 = _GEN_1545[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1546 = {1{$random}};
  inputMemBlock_7 = _GEN_1546[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1547 = {1{$random}};
  inputMemBlock_8 = _GEN_1547[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1548 = {1{$random}};
  inputMemBlock_9 = _GEN_1548[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1549 = {1{$random}};
  inputMemBlock_10 = _GEN_1549[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1550 = {1{$random}};
  inputMemBlock_11 = _GEN_1550[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1551 = {1{$random}};
  inputMemBlock_12 = _GEN_1551[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1552 = {1{$random}};
  inputMemBlock_13 = _GEN_1552[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1553 = {1{$random}};
  inputMemBlock_14 = _GEN_1553[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1554 = {1{$random}};
  inputMemBlock_15 = _GEN_1554[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1555 = {1{$random}};
  inputMemBlock_16 = _GEN_1555[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1556 = {1{$random}};
  inputMemBlock_17 = _GEN_1556[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1557 = {1{$random}};
  inputMemBlock_18 = _GEN_1557[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1558 = {1{$random}};
  inputMemBlock_19 = _GEN_1558[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1559 = {1{$random}};
  inputMemBlock_20 = _GEN_1559[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1560 = {1{$random}};
  inputMemBlock_21 = _GEN_1560[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1561 = {1{$random}};
  inputMemBlock_22 = _GEN_1561[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1562 = {1{$random}};
  inputMemBlock_23 = _GEN_1562[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1563 = {1{$random}};
  inputMemBlock_24 = _GEN_1563[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1564 = {1{$random}};
  inputMemBlock_25 = _GEN_1564[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1565 = {1{$random}};
  inputMemBlock_26 = _GEN_1565[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1566 = {1{$random}};
  inputMemBlock_27 = _GEN_1566[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1567 = {1{$random}};
  inputMemBlock_28 = _GEN_1567[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1568 = {1{$random}};
  inputMemBlock_29 = _GEN_1568[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1569 = {1{$random}};
  inputMemBlock_30 = _GEN_1569[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1570 = {1{$random}};
  inputMemBlock_31 = _GEN_1570[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1571 = {1{$random}};
  inputMemBlock_32 = _GEN_1571[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1572 = {1{$random}};
  inputMemBlock_33 = _GEN_1572[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1573 = {1{$random}};
  inputMemBlock_34 = _GEN_1573[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1574 = {1{$random}};
  inputMemBlock_35 = _GEN_1574[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1575 = {1{$random}};
  inputMemBlock_36 = _GEN_1575[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1576 = {1{$random}};
  inputMemBlock_37 = _GEN_1576[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1577 = {1{$random}};
  inputMemBlock_38 = _GEN_1577[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1578 = {1{$random}};
  inputMemBlock_39 = _GEN_1578[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1579 = {1{$random}};
  inputMemBlock_40 = _GEN_1579[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1580 = {1{$random}};
  inputMemBlock_41 = _GEN_1580[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1581 = {1{$random}};
  inputMemBlock_42 = _GEN_1581[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1582 = {1{$random}};
  inputMemBlock_43 = _GEN_1582[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1583 = {1{$random}};
  inputMemBlock_44 = _GEN_1583[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1584 = {1{$random}};
  inputMemBlock_45 = _GEN_1584[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1585 = {1{$random}};
  inputMemBlock_46 = _GEN_1585[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1586 = {1{$random}};
  inputMemBlock_47 = _GEN_1586[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1587 = {1{$random}};
  inputMemBlock_48 = _GEN_1587[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1588 = {1{$random}};
  inputMemBlock_49 = _GEN_1588[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1589 = {1{$random}};
  inputMemBlock_50 = _GEN_1589[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1590 = {1{$random}};
  inputMemBlock_51 = _GEN_1590[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1591 = {1{$random}};
  inputMemBlock_52 = _GEN_1591[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1592 = {1{$random}};
  inputMemBlock_53 = _GEN_1592[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1593 = {1{$random}};
  inputMemBlock_54 = _GEN_1593[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1594 = {1{$random}};
  inputMemBlock_55 = _GEN_1594[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1595 = {1{$random}};
  inputMemBlock_56 = _GEN_1595[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1596 = {1{$random}};
  inputMemBlock_57 = _GEN_1596[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1597 = {1{$random}};
  inputMemBlock_58 = _GEN_1597[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1598 = {1{$random}};
  inputMemBlock_59 = _GEN_1598[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1599 = {1{$random}};
  inputMemBlock_60 = _GEN_1599[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1600 = {1{$random}};
  inputMemBlock_61 = _GEN_1600[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1601 = {1{$random}};
  inputMemBlock_62 = _GEN_1601[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1602 = {1{$random}};
  inputMemBlock_63 = _GEN_1602[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1603 = {1{$random}};
  inputMemBlock_64 = _GEN_1603[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1604 = {1{$random}};
  inputMemBlock_65 = _GEN_1604[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1605 = {1{$random}};
  inputMemBlock_66 = _GEN_1605[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1606 = {1{$random}};
  inputMemBlock_67 = _GEN_1606[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1607 = {1{$random}};
  inputMemBlock_68 = _GEN_1607[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1608 = {1{$random}};
  inputMemBlock_69 = _GEN_1608[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1609 = {1{$random}};
  inputMemBlock_70 = _GEN_1609[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1610 = {1{$random}};
  inputMemBlock_71 = _GEN_1610[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1611 = {1{$random}};
  inputMemBlock_72 = _GEN_1611[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1612 = {1{$random}};
  inputMemBlock_73 = _GEN_1612[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1613 = {1{$random}};
  inputMemBlock_74 = _GEN_1613[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1614 = {1{$random}};
  inputMemBlock_75 = _GEN_1614[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1615 = {1{$random}};
  inputMemBlock_76 = _GEN_1615[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1616 = {1{$random}};
  inputMemBlock_77 = _GEN_1616[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1617 = {1{$random}};
  inputMemBlock_78 = _GEN_1617[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1618 = {1{$random}};
  inputMemBlock_79 = _GEN_1618[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1619 = {1{$random}};
  inputMemBlock_80 = _GEN_1619[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1620 = {1{$random}};
  inputMemBlock_81 = _GEN_1620[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1621 = {1{$random}};
  inputMemBlock_82 = _GEN_1621[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1622 = {1{$random}};
  inputMemBlock_83 = _GEN_1622[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1623 = {1{$random}};
  inputMemBlock_84 = _GEN_1623[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1624 = {1{$random}};
  inputMemBlock_85 = _GEN_1624[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1625 = {1{$random}};
  inputMemBlock_86 = _GEN_1625[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1626 = {1{$random}};
  inputMemBlock_87 = _GEN_1626[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1627 = {1{$random}};
  inputMemBlock_88 = _GEN_1627[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1628 = {1{$random}};
  inputMemBlock_89 = _GEN_1628[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1629 = {1{$random}};
  inputMemBlock_90 = _GEN_1629[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1630 = {1{$random}};
  inputMemBlock_91 = _GEN_1630[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1631 = {1{$random}};
  inputMemBlock_92 = _GEN_1631[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1632 = {1{$random}};
  inputMemBlock_93 = _GEN_1632[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1633 = {1{$random}};
  inputMemBlock_94 = _GEN_1633[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1634 = {1{$random}};
  inputMemBlock_95 = _GEN_1634[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1635 = {1{$random}};
  inputMemBlock_96 = _GEN_1635[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1636 = {1{$random}};
  inputMemBlock_97 = _GEN_1636[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1637 = {1{$random}};
  inputMemBlock_98 = _GEN_1637[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1638 = {1{$random}};
  inputMemBlock_99 = _GEN_1638[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1639 = {1{$random}};
  inputMemBlock_100 = _GEN_1639[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1640 = {1{$random}};
  inputMemBlock_101 = _GEN_1640[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1641 = {1{$random}};
  inputMemBlock_102 = _GEN_1641[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1642 = {1{$random}};
  inputMemBlock_103 = _GEN_1642[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1643 = {1{$random}};
  inputMemBlock_104 = _GEN_1643[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1644 = {1{$random}};
  inputMemBlock_105 = _GEN_1644[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1645 = {1{$random}};
  inputMemBlock_106 = _GEN_1645[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1646 = {1{$random}};
  inputMemBlock_107 = _GEN_1646[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1647 = {1{$random}};
  inputMemBlock_108 = _GEN_1647[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1648 = {1{$random}};
  inputMemBlock_109 = _GEN_1648[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1649 = {1{$random}};
  inputMemBlock_110 = _GEN_1649[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1650 = {1{$random}};
  inputMemBlock_111 = _GEN_1650[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1651 = {1{$random}};
  inputMemBlock_112 = _GEN_1651[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1652 = {1{$random}};
  inputMemBlock_113 = _GEN_1652[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1653 = {1{$random}};
  inputMemBlock_114 = _GEN_1653[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1654 = {1{$random}};
  inputMemBlock_115 = _GEN_1654[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1655 = {1{$random}};
  inputMemBlock_116 = _GEN_1655[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1656 = {1{$random}};
  inputMemBlock_117 = _GEN_1656[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1657 = {1{$random}};
  inputMemBlock_118 = _GEN_1657[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1658 = {1{$random}};
  inputMemBlock_119 = _GEN_1658[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1659 = {1{$random}};
  inputMemBlock_120 = _GEN_1659[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1660 = {1{$random}};
  inputMemBlock_121 = _GEN_1660[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1661 = {1{$random}};
  inputMemBlock_122 = _GEN_1661[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1662 = {1{$random}};
  inputMemBlock_123 = _GEN_1662[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1663 = {1{$random}};
  inputMemBlock_124 = _GEN_1663[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1664 = {1{$random}};
  inputMemBlock_125 = _GEN_1664[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1665 = {1{$random}};
  inputMemBlock_126 = _GEN_1665[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1666 = {1{$random}};
  inputMemBlock_127 = _GEN_1666[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1667 = {1{$random}};
  inputMemBlock_128 = _GEN_1667[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1668 = {1{$random}};
  inputMemBlock_129 = _GEN_1668[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1669 = {1{$random}};
  inputMemBlock_130 = _GEN_1669[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1670 = {1{$random}};
  inputMemBlock_131 = _GEN_1670[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1671 = {1{$random}};
  inputMemBlock_132 = _GEN_1671[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1672 = {1{$random}};
  inputMemBlock_133 = _GEN_1672[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1673 = {1{$random}};
  inputMemBlock_134 = _GEN_1673[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1674 = {1{$random}};
  inputMemBlock_135 = _GEN_1674[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1675 = {1{$random}};
  inputMemBlock_136 = _GEN_1675[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1676 = {1{$random}};
  inputMemBlock_137 = _GEN_1676[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1677 = {1{$random}};
  inputMemBlock_138 = _GEN_1677[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1678 = {1{$random}};
  inputMemBlock_139 = _GEN_1678[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1679 = {1{$random}};
  inputMemBlock_140 = _GEN_1679[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1680 = {1{$random}};
  inputMemBlock_141 = _GEN_1680[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1681 = {1{$random}};
  inputMemBlock_142 = _GEN_1681[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1682 = {1{$random}};
  inputMemBlock_143 = _GEN_1682[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1683 = {1{$random}};
  inputMemBlock_144 = _GEN_1683[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1684 = {1{$random}};
  inputMemBlock_145 = _GEN_1684[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1685 = {1{$random}};
  inputMemBlock_146 = _GEN_1685[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1686 = {1{$random}};
  inputMemBlock_147 = _GEN_1686[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1687 = {1{$random}};
  inputMemBlock_148 = _GEN_1687[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1688 = {1{$random}};
  inputMemBlock_149 = _GEN_1688[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1689 = {1{$random}};
  inputMemBlock_150 = _GEN_1689[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1690 = {1{$random}};
  inputMemBlock_151 = _GEN_1690[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1691 = {1{$random}};
  inputMemBlock_152 = _GEN_1691[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1692 = {1{$random}};
  inputMemBlock_153 = _GEN_1692[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1693 = {1{$random}};
  inputMemBlock_154 = _GEN_1693[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1694 = {1{$random}};
  inputMemBlock_155 = _GEN_1694[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1695 = {1{$random}};
  inputMemBlock_156 = _GEN_1695[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1696 = {1{$random}};
  inputMemBlock_157 = _GEN_1696[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1697 = {1{$random}};
  inputMemBlock_158 = _GEN_1697[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1698 = {1{$random}};
  inputMemBlock_159 = _GEN_1698[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1699 = {1{$random}};
  inputMemBlock_160 = _GEN_1699[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1700 = {1{$random}};
  inputMemBlock_161 = _GEN_1700[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1701 = {1{$random}};
  inputMemBlock_162 = _GEN_1701[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1702 = {1{$random}};
  inputMemBlock_163 = _GEN_1702[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1703 = {1{$random}};
  inputMemBlock_164 = _GEN_1703[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1704 = {1{$random}};
  inputMemBlock_165 = _GEN_1704[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1705 = {1{$random}};
  inputMemBlock_166 = _GEN_1705[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1706 = {1{$random}};
  inputMemBlock_167 = _GEN_1706[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1707 = {1{$random}};
  inputMemBlock_168 = _GEN_1707[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1708 = {1{$random}};
  inputMemBlock_169 = _GEN_1708[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1709 = {1{$random}};
  inputMemBlock_170 = _GEN_1709[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1710 = {1{$random}};
  inputMemBlock_171 = _GEN_1710[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1711 = {1{$random}};
  inputMemBlock_172 = _GEN_1711[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1712 = {1{$random}};
  inputMemBlock_173 = _GEN_1712[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1713 = {1{$random}};
  inputMemBlock_174 = _GEN_1713[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1714 = {1{$random}};
  inputMemBlock_175 = _GEN_1714[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1715 = {1{$random}};
  inputMemBlock_176 = _GEN_1715[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1716 = {1{$random}};
  inputMemBlock_177 = _GEN_1716[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1717 = {1{$random}};
  inputMemBlock_178 = _GEN_1717[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1718 = {1{$random}};
  inputMemBlock_179 = _GEN_1718[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1719 = {1{$random}};
  inputMemBlock_180 = _GEN_1719[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1720 = {1{$random}};
  inputMemBlock_181 = _GEN_1720[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1721 = {1{$random}};
  inputMemBlock_182 = _GEN_1721[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1722 = {1{$random}};
  inputMemBlock_183 = _GEN_1722[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1723 = {1{$random}};
  inputMemBlock_184 = _GEN_1723[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1724 = {1{$random}};
  inputMemBlock_185 = _GEN_1724[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1725 = {1{$random}};
  inputMemBlock_186 = _GEN_1725[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1726 = {1{$random}};
  inputMemBlock_187 = _GEN_1726[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1727 = {1{$random}};
  inputMemBlock_188 = _GEN_1727[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1728 = {1{$random}};
  inputMemBlock_189 = _GEN_1728[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1729 = {1{$random}};
  inputMemBlock_190 = _GEN_1729[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1730 = {1{$random}};
  inputMemBlock_191 = _GEN_1730[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1731 = {1{$random}};
  inputMemBlock_192 = _GEN_1731[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1732 = {1{$random}};
  inputMemBlock_193 = _GEN_1732[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1733 = {1{$random}};
  inputMemBlock_194 = _GEN_1733[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1734 = {1{$random}};
  inputMemBlock_195 = _GEN_1734[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1735 = {1{$random}};
  inputMemBlock_196 = _GEN_1735[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1736 = {1{$random}};
  inputMemBlock_197 = _GEN_1736[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1737 = {1{$random}};
  inputMemBlock_198 = _GEN_1737[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1738 = {1{$random}};
  inputMemBlock_199 = _GEN_1738[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1739 = {1{$random}};
  inputMemBlock_200 = _GEN_1739[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1740 = {1{$random}};
  inputMemBlock_201 = _GEN_1740[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1741 = {1{$random}};
  inputMemBlock_202 = _GEN_1741[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1742 = {1{$random}};
  inputMemBlock_203 = _GEN_1742[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1743 = {1{$random}};
  inputMemBlock_204 = _GEN_1743[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1744 = {1{$random}};
  inputMemBlock_205 = _GEN_1744[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1745 = {1{$random}};
  inputMemBlock_206 = _GEN_1745[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1746 = {1{$random}};
  inputMemBlock_207 = _GEN_1746[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1747 = {1{$random}};
  inputMemBlock_208 = _GEN_1747[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1748 = {1{$random}};
  inputMemBlock_209 = _GEN_1748[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1749 = {1{$random}};
  inputMemBlock_210 = _GEN_1749[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1750 = {1{$random}};
  inputMemBlock_211 = _GEN_1750[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1751 = {1{$random}};
  inputMemBlock_212 = _GEN_1751[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1752 = {1{$random}};
  inputMemBlock_213 = _GEN_1752[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1753 = {1{$random}};
  inputMemBlock_214 = _GEN_1753[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1754 = {1{$random}};
  inputMemBlock_215 = _GEN_1754[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1755 = {1{$random}};
  inputMemBlock_216 = _GEN_1755[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1756 = {1{$random}};
  inputMemBlock_217 = _GEN_1756[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1757 = {1{$random}};
  inputMemBlock_218 = _GEN_1757[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1758 = {1{$random}};
  inputMemBlock_219 = _GEN_1758[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1759 = {1{$random}};
  inputMemBlock_220 = _GEN_1759[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1760 = {1{$random}};
  inputMemBlock_221 = _GEN_1760[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1761 = {1{$random}};
  inputMemBlock_222 = _GEN_1761[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1762 = {1{$random}};
  inputMemBlock_223 = _GEN_1762[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1763 = {1{$random}};
  inputMemBlock_224 = _GEN_1763[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1764 = {1{$random}};
  inputMemBlock_225 = _GEN_1764[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1765 = {1{$random}};
  inputMemBlock_226 = _GEN_1765[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1766 = {1{$random}};
  inputMemBlock_227 = _GEN_1766[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1767 = {1{$random}};
  inputMemBlock_228 = _GEN_1767[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1768 = {1{$random}};
  inputMemBlock_229 = _GEN_1768[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1769 = {1{$random}};
  inputMemBlock_230 = _GEN_1769[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1770 = {1{$random}};
  inputMemBlock_231 = _GEN_1770[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1771 = {1{$random}};
  inputMemBlock_232 = _GEN_1771[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1772 = {1{$random}};
  inputMemBlock_233 = _GEN_1772[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1773 = {1{$random}};
  inputMemBlock_234 = _GEN_1773[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1774 = {1{$random}};
  inputMemBlock_235 = _GEN_1774[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1775 = {1{$random}};
  inputMemBlock_236 = _GEN_1775[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1776 = {1{$random}};
  inputMemBlock_237 = _GEN_1776[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1777 = {1{$random}};
  inputMemBlock_238 = _GEN_1777[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1778 = {1{$random}};
  inputMemBlock_239 = _GEN_1778[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1779 = {1{$random}};
  inputMemBlock_240 = _GEN_1779[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1780 = {1{$random}};
  inputMemBlock_241 = _GEN_1780[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1781 = {1{$random}};
  inputMemBlock_242 = _GEN_1781[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1782 = {1{$random}};
  inputMemBlock_243 = _GEN_1782[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1783 = {1{$random}};
  inputMemBlock_244 = _GEN_1783[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1784 = {1{$random}};
  inputMemBlock_245 = _GEN_1784[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1785 = {1{$random}};
  inputMemBlock_246 = _GEN_1785[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1786 = {1{$random}};
  inputMemBlock_247 = _GEN_1786[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1787 = {1{$random}};
  inputMemBlock_248 = _GEN_1787[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1788 = {1{$random}};
  inputMemBlock_249 = _GEN_1788[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1789 = {1{$random}};
  inputMemBlock_250 = _GEN_1789[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1790 = {1{$random}};
  inputMemBlock_251 = _GEN_1790[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1791 = {1{$random}};
  inputMemBlock_252 = _GEN_1791[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1792 = {1{$random}};
  inputMemBlock_253 = _GEN_1792[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1793 = {1{$random}};
  inputMemBlock_254 = _GEN_1793[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1794 = {1{$random}};
  inputMemBlock_255 = _GEN_1794[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1795 = {1{$random}};
  inputMemBlock_256 = _GEN_1795[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1796 = {1{$random}};
  inputMemBlock_257 = _GEN_1796[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1797 = {1{$random}};
  inputMemBlock_258 = _GEN_1797[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1798 = {1{$random}};
  inputMemBlock_259 = _GEN_1798[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1799 = {1{$random}};
  inputMemBlock_260 = _GEN_1799[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1800 = {1{$random}};
  inputMemBlock_261 = _GEN_1800[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1801 = {1{$random}};
  inputMemBlock_262 = _GEN_1801[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1802 = {1{$random}};
  inputMemBlock_263 = _GEN_1802[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1803 = {1{$random}};
  inputMemBlock_264 = _GEN_1803[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1804 = {1{$random}};
  inputMemBlock_265 = _GEN_1804[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1805 = {1{$random}};
  inputMemBlock_266 = _GEN_1805[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1806 = {1{$random}};
  inputMemBlock_267 = _GEN_1806[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1807 = {1{$random}};
  inputMemBlock_268 = _GEN_1807[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1808 = {1{$random}};
  inputMemBlock_269 = _GEN_1808[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1809 = {1{$random}};
  inputMemBlock_270 = _GEN_1809[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1810 = {1{$random}};
  inputMemBlock_271 = _GEN_1810[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1811 = {1{$random}};
  inputMemBlock_272 = _GEN_1811[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1812 = {1{$random}};
  inputMemBlock_273 = _GEN_1812[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1813 = {1{$random}};
  inputMemBlock_274 = _GEN_1813[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1814 = {1{$random}};
  inputMemBlock_275 = _GEN_1814[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1815 = {1{$random}};
  inputMemBlock_276 = _GEN_1815[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1816 = {1{$random}};
  inputMemBlock_277 = _GEN_1816[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1817 = {1{$random}};
  inputMemBlock_278 = _GEN_1817[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1818 = {1{$random}};
  inputMemBlock_279 = _GEN_1818[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1819 = {1{$random}};
  inputMemBlock_280 = _GEN_1819[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1820 = {1{$random}};
  inputMemBlock_281 = _GEN_1820[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1821 = {1{$random}};
  inputMemBlock_282 = _GEN_1821[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1822 = {1{$random}};
  inputMemBlock_283 = _GEN_1822[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1823 = {1{$random}};
  inputMemBlock_284 = _GEN_1823[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1824 = {1{$random}};
  inputMemBlock_285 = _GEN_1824[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1825 = {1{$random}};
  inputMemBlock_286 = _GEN_1825[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1826 = {1{$random}};
  inputMemBlock_287 = _GEN_1826[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1827 = {1{$random}};
  inputMemBlock_288 = _GEN_1827[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1828 = {1{$random}};
  inputMemBlock_289 = _GEN_1828[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1829 = {1{$random}};
  inputMemBlock_290 = _GEN_1829[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1830 = {1{$random}};
  inputMemBlock_291 = _GEN_1830[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1831 = {1{$random}};
  inputMemBlock_292 = _GEN_1831[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1832 = {1{$random}};
  inputMemBlock_293 = _GEN_1832[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1833 = {1{$random}};
  inputMemBlock_294 = _GEN_1833[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1834 = {1{$random}};
  inputMemBlock_295 = _GEN_1834[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1835 = {1{$random}};
  inputMemBlock_296 = _GEN_1835[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1836 = {1{$random}};
  inputMemBlock_297 = _GEN_1836[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1837 = {1{$random}};
  inputMemBlock_298 = _GEN_1837[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1838 = {1{$random}};
  inputMemBlock_299 = _GEN_1838[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1839 = {1{$random}};
  inputMemBlock_300 = _GEN_1839[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1840 = {1{$random}};
  inputMemBlock_301 = _GEN_1840[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1841 = {1{$random}};
  inputMemBlock_302 = _GEN_1841[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1842 = {1{$random}};
  inputMemBlock_303 = _GEN_1842[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1843 = {1{$random}};
  inputMemBlock_304 = _GEN_1843[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1844 = {1{$random}};
  inputMemBlock_305 = _GEN_1844[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1845 = {1{$random}};
  inputMemBlock_306 = _GEN_1845[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1846 = {1{$random}};
  inputMemBlock_307 = _GEN_1846[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1847 = {1{$random}};
  inputMemBlock_308 = _GEN_1847[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1848 = {1{$random}};
  inputMemBlock_309 = _GEN_1848[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1849 = {1{$random}};
  inputMemBlock_310 = _GEN_1849[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1850 = {1{$random}};
  inputMemBlock_311 = _GEN_1850[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1851 = {1{$random}};
  inputMemBlock_312 = _GEN_1851[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1852 = {1{$random}};
  inputMemBlock_313 = _GEN_1852[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1853 = {1{$random}};
  inputMemBlock_314 = _GEN_1853[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1854 = {1{$random}};
  inputMemBlock_315 = _GEN_1854[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1855 = {1{$random}};
  inputMemBlock_316 = _GEN_1855[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1856 = {1{$random}};
  inputMemBlock_317 = _GEN_1856[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1857 = {1{$random}};
  inputMemBlock_318 = _GEN_1857[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1858 = {1{$random}};
  inputMemBlock_319 = _GEN_1858[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1859 = {1{$random}};
  inputMemBlock_320 = _GEN_1859[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1860 = {1{$random}};
  inputMemBlock_321 = _GEN_1860[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1861 = {1{$random}};
  inputMemBlock_322 = _GEN_1861[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1862 = {1{$random}};
  inputMemBlock_323 = _GEN_1862[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1863 = {1{$random}};
  inputMemBlock_324 = _GEN_1863[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1864 = {1{$random}};
  inputMemBlock_325 = _GEN_1864[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1865 = {1{$random}};
  inputMemBlock_326 = _GEN_1865[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1866 = {1{$random}};
  inputMemBlock_327 = _GEN_1866[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1867 = {1{$random}};
  inputMemBlock_328 = _GEN_1867[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1868 = {1{$random}};
  inputMemBlock_329 = _GEN_1868[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1869 = {1{$random}};
  inputMemBlock_330 = _GEN_1869[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1870 = {1{$random}};
  inputMemBlock_331 = _GEN_1870[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1871 = {1{$random}};
  inputMemBlock_332 = _GEN_1871[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1872 = {1{$random}};
  inputMemBlock_333 = _GEN_1872[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1873 = {1{$random}};
  inputMemBlock_334 = _GEN_1873[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1874 = {1{$random}};
  inputMemBlock_335 = _GEN_1874[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1875 = {1{$random}};
  inputMemBlock_336 = _GEN_1875[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1876 = {1{$random}};
  inputMemBlock_337 = _GEN_1876[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1877 = {1{$random}};
  inputMemBlock_338 = _GEN_1877[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1878 = {1{$random}};
  inputMemBlock_339 = _GEN_1878[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1879 = {1{$random}};
  inputMemBlock_340 = _GEN_1879[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1880 = {1{$random}};
  inputMemBlock_341 = _GEN_1880[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1881 = {1{$random}};
  inputMemBlock_342 = _GEN_1881[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1882 = {1{$random}};
  inputMemBlock_343 = _GEN_1882[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1883 = {1{$random}};
  inputMemBlock_344 = _GEN_1883[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1884 = {1{$random}};
  inputMemBlock_345 = _GEN_1884[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1885 = {1{$random}};
  inputMemBlock_346 = _GEN_1885[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1886 = {1{$random}};
  inputMemBlock_347 = _GEN_1886[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1887 = {1{$random}};
  inputMemBlock_348 = _GEN_1887[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1888 = {1{$random}};
  inputMemBlock_349 = _GEN_1888[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1889 = {1{$random}};
  inputMemBlock_350 = _GEN_1889[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1890 = {1{$random}};
  inputMemBlock_351 = _GEN_1890[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1891 = {1{$random}};
  inputMemBlock_352 = _GEN_1891[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1892 = {1{$random}};
  inputMemBlock_353 = _GEN_1892[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1893 = {1{$random}};
  inputMemBlock_354 = _GEN_1893[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1894 = {1{$random}};
  inputMemBlock_355 = _GEN_1894[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1895 = {1{$random}};
  inputMemBlock_356 = _GEN_1895[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1896 = {1{$random}};
  inputMemBlock_357 = _GEN_1896[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1897 = {1{$random}};
  inputMemBlock_358 = _GEN_1897[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1898 = {1{$random}};
  inputMemBlock_359 = _GEN_1898[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1899 = {1{$random}};
  inputMemBlock_360 = _GEN_1899[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1900 = {1{$random}};
  inputMemBlock_361 = _GEN_1900[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1901 = {1{$random}};
  inputMemBlock_362 = _GEN_1901[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1902 = {1{$random}};
  inputMemBlock_363 = _GEN_1902[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1903 = {1{$random}};
  inputMemBlock_364 = _GEN_1903[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1904 = {1{$random}};
  inputMemBlock_365 = _GEN_1904[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1905 = {1{$random}};
  inputMemBlock_366 = _GEN_1905[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1906 = {1{$random}};
  inputMemBlock_367 = _GEN_1906[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1907 = {1{$random}};
  inputMemBlock_368 = _GEN_1907[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1908 = {1{$random}};
  inputMemBlock_369 = _GEN_1908[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1909 = {1{$random}};
  inputMemBlock_370 = _GEN_1909[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1910 = {1{$random}};
  inputMemBlock_371 = _GEN_1910[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1911 = {1{$random}};
  inputMemBlock_372 = _GEN_1911[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1912 = {1{$random}};
  inputMemBlock_373 = _GEN_1912[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1913 = {1{$random}};
  inputMemBlock_374 = _GEN_1913[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1914 = {1{$random}};
  inputMemBlock_375 = _GEN_1914[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1915 = {1{$random}};
  inputMemBlock_376 = _GEN_1915[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1916 = {1{$random}};
  inputMemBlock_377 = _GEN_1916[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1917 = {1{$random}};
  inputMemBlock_378 = _GEN_1917[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1918 = {1{$random}};
  inputMemBlock_379 = _GEN_1918[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1919 = {1{$random}};
  inputMemBlock_380 = _GEN_1919[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1920 = {1{$random}};
  inputMemBlock_381 = _GEN_1920[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1921 = {1{$random}};
  inputMemBlock_382 = _GEN_1921[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1922 = {1{$random}};
  inputMemBlock_383 = _GEN_1922[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1923 = {1{$random}};
  inputMemBlock_384 = _GEN_1923[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1924 = {1{$random}};
  inputMemBlock_385 = _GEN_1924[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1925 = {1{$random}};
  inputMemBlock_386 = _GEN_1925[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1926 = {1{$random}};
  inputMemBlock_387 = _GEN_1926[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1927 = {1{$random}};
  inputMemBlock_388 = _GEN_1927[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1928 = {1{$random}};
  inputMemBlock_389 = _GEN_1928[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1929 = {1{$random}};
  inputMemBlock_390 = _GEN_1929[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1930 = {1{$random}};
  inputMemBlock_391 = _GEN_1930[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1931 = {1{$random}};
  inputMemBlock_392 = _GEN_1931[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1932 = {1{$random}};
  inputMemBlock_393 = _GEN_1932[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1933 = {1{$random}};
  inputMemBlock_394 = _GEN_1933[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1934 = {1{$random}};
  inputMemBlock_395 = _GEN_1934[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1935 = {1{$random}};
  inputMemBlock_396 = _GEN_1935[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1936 = {1{$random}};
  inputMemBlock_397 = _GEN_1936[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1937 = {1{$random}};
  inputMemBlock_398 = _GEN_1937[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1938 = {1{$random}};
  inputMemBlock_399 = _GEN_1938[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1939 = {1{$random}};
  inputMemBlock_400 = _GEN_1939[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1940 = {1{$random}};
  inputMemBlock_401 = _GEN_1940[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1941 = {1{$random}};
  inputMemBlock_402 = _GEN_1941[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1942 = {1{$random}};
  inputMemBlock_403 = _GEN_1942[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1943 = {1{$random}};
  inputMemBlock_404 = _GEN_1943[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1944 = {1{$random}};
  inputMemBlock_405 = _GEN_1944[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1945 = {1{$random}};
  inputMemBlock_406 = _GEN_1945[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1946 = {1{$random}};
  inputMemBlock_407 = _GEN_1946[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1947 = {1{$random}};
  inputMemBlock_408 = _GEN_1947[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1948 = {1{$random}};
  inputMemBlock_409 = _GEN_1948[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1949 = {1{$random}};
  inputMemBlock_410 = _GEN_1949[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1950 = {1{$random}};
  inputMemBlock_411 = _GEN_1950[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1951 = {1{$random}};
  inputMemBlock_412 = _GEN_1951[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1952 = {1{$random}};
  inputMemBlock_413 = _GEN_1952[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1953 = {1{$random}};
  inputMemBlock_414 = _GEN_1953[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1954 = {1{$random}};
  inputMemBlock_415 = _GEN_1954[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1955 = {1{$random}};
  inputMemBlock_416 = _GEN_1955[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1956 = {1{$random}};
  inputMemBlock_417 = _GEN_1956[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1957 = {1{$random}};
  inputMemBlock_418 = _GEN_1957[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1958 = {1{$random}};
  inputMemBlock_419 = _GEN_1958[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1959 = {1{$random}};
  inputMemBlock_420 = _GEN_1959[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1960 = {1{$random}};
  inputMemBlock_421 = _GEN_1960[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1961 = {1{$random}};
  inputMemBlock_422 = _GEN_1961[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1962 = {1{$random}};
  inputMemBlock_423 = _GEN_1962[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1963 = {1{$random}};
  inputMemBlock_424 = _GEN_1963[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1964 = {1{$random}};
  inputMemBlock_425 = _GEN_1964[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1965 = {1{$random}};
  inputMemBlock_426 = _GEN_1965[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1966 = {1{$random}};
  inputMemBlock_427 = _GEN_1966[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1967 = {1{$random}};
  inputMemBlock_428 = _GEN_1967[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1968 = {1{$random}};
  inputMemBlock_429 = _GEN_1968[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1969 = {1{$random}};
  inputMemBlock_430 = _GEN_1969[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1970 = {1{$random}};
  inputMemBlock_431 = _GEN_1970[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1971 = {1{$random}};
  inputMemBlock_432 = _GEN_1971[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1972 = {1{$random}};
  inputMemBlock_433 = _GEN_1972[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1973 = {1{$random}};
  inputMemBlock_434 = _GEN_1973[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1974 = {1{$random}};
  inputMemBlock_435 = _GEN_1974[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1975 = {1{$random}};
  inputMemBlock_436 = _GEN_1975[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1976 = {1{$random}};
  inputMemBlock_437 = _GEN_1976[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1977 = {1{$random}};
  inputMemBlock_438 = _GEN_1977[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1978 = {1{$random}};
  inputMemBlock_439 = _GEN_1978[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1979 = {1{$random}};
  inputMemBlock_440 = _GEN_1979[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1980 = {1{$random}};
  inputMemBlock_441 = _GEN_1980[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1981 = {1{$random}};
  inputMemBlock_442 = _GEN_1981[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1982 = {1{$random}};
  inputMemBlock_443 = _GEN_1982[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1983 = {1{$random}};
  inputMemBlock_444 = _GEN_1983[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1984 = {1{$random}};
  inputMemBlock_445 = _GEN_1984[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1985 = {1{$random}};
  inputMemBlock_446 = _GEN_1985[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1986 = {1{$random}};
  inputMemBlock_447 = _GEN_1986[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1987 = {1{$random}};
  inputMemBlock_448 = _GEN_1987[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1988 = {1{$random}};
  inputMemBlock_449 = _GEN_1988[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1989 = {1{$random}};
  inputMemBlock_450 = _GEN_1989[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1990 = {1{$random}};
  inputMemBlock_451 = _GEN_1990[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1991 = {1{$random}};
  inputMemBlock_452 = _GEN_1991[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1992 = {1{$random}};
  inputMemBlock_453 = _GEN_1992[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1993 = {1{$random}};
  inputMemBlock_454 = _GEN_1993[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1994 = {1{$random}};
  inputMemBlock_455 = _GEN_1994[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1995 = {1{$random}};
  inputMemBlock_456 = _GEN_1995[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1996 = {1{$random}};
  inputMemBlock_457 = _GEN_1996[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1997 = {1{$random}};
  inputMemBlock_458 = _GEN_1997[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1998 = {1{$random}};
  inputMemBlock_459 = _GEN_1998[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1999 = {1{$random}};
  inputMemBlock_460 = _GEN_1999[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2000 = {1{$random}};
  inputMemBlock_461 = _GEN_2000[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2001 = {1{$random}};
  inputMemBlock_462 = _GEN_2001[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2002 = {1{$random}};
  inputMemBlock_463 = _GEN_2002[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2003 = {1{$random}};
  inputMemBlock_464 = _GEN_2003[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2004 = {1{$random}};
  inputMemBlock_465 = _GEN_2004[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2005 = {1{$random}};
  inputMemBlock_466 = _GEN_2005[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2006 = {1{$random}};
  inputMemBlock_467 = _GEN_2006[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2007 = {1{$random}};
  inputMemBlock_468 = _GEN_2007[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2008 = {1{$random}};
  inputMemBlock_469 = _GEN_2008[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2009 = {1{$random}};
  inputMemBlock_470 = _GEN_2009[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2010 = {1{$random}};
  inputMemBlock_471 = _GEN_2010[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2011 = {1{$random}};
  inputMemBlock_472 = _GEN_2011[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2012 = {1{$random}};
  inputMemBlock_473 = _GEN_2012[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2013 = {1{$random}};
  inputMemBlock_474 = _GEN_2013[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2014 = {1{$random}};
  inputMemBlock_475 = _GEN_2014[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2015 = {1{$random}};
  inputMemBlock_476 = _GEN_2015[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2016 = {1{$random}};
  inputMemBlock_477 = _GEN_2016[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2017 = {1{$random}};
  inputMemBlock_478 = _GEN_2017[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2018 = {1{$random}};
  inputMemBlock_479 = _GEN_2018[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2019 = {1{$random}};
  inputMemBlock_480 = _GEN_2019[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2020 = {1{$random}};
  inputMemBlock_481 = _GEN_2020[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2021 = {1{$random}};
  inputMemBlock_482 = _GEN_2021[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2022 = {1{$random}};
  inputMemBlock_483 = _GEN_2022[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2023 = {1{$random}};
  inputMemBlock_484 = _GEN_2023[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2024 = {1{$random}};
  inputMemBlock_485 = _GEN_2024[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2025 = {1{$random}};
  inputMemBlock_486 = _GEN_2025[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2026 = {1{$random}};
  inputMemBlock_487 = _GEN_2026[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2027 = {1{$random}};
  inputMemBlock_488 = _GEN_2027[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2028 = {1{$random}};
  inputMemBlock_489 = _GEN_2028[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2029 = {1{$random}};
  inputMemBlock_490 = _GEN_2029[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2030 = {1{$random}};
  inputMemBlock_491 = _GEN_2030[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2031 = {1{$random}};
  inputMemBlock_492 = _GEN_2031[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2032 = {1{$random}};
  inputMemBlock_493 = _GEN_2032[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2033 = {1{$random}};
  inputMemBlock_494 = _GEN_2033[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2034 = {1{$random}};
  inputMemBlock_495 = _GEN_2034[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2035 = {1{$random}};
  inputMemBlock_496 = _GEN_2035[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2036 = {1{$random}};
  inputMemBlock_497 = _GEN_2036[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2037 = {1{$random}};
  inputMemBlock_498 = _GEN_2037[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2038 = {1{$random}};
  inputMemBlock_499 = _GEN_2038[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2039 = {1{$random}};
  inputMemBlock_500 = _GEN_2039[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2040 = {1{$random}};
  inputMemBlock_501 = _GEN_2040[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2041 = {1{$random}};
  inputMemBlock_502 = _GEN_2041[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2042 = {1{$random}};
  inputMemBlock_503 = _GEN_2042[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2043 = {1{$random}};
  inputMemBlock_504 = _GEN_2043[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2044 = {1{$random}};
  inputMemBlock_505 = _GEN_2044[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2045 = {1{$random}};
  inputMemBlock_506 = _GEN_2045[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2046 = {1{$random}};
  inputMemBlock_507 = _GEN_2046[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2047 = {1{$random}};
  inputMemBlock_508 = _GEN_2047[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2048 = {1{$random}};
  inputMemBlock_509 = _GEN_2048[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2049 = {1{$random}};
  inputMemBlock_510 = _GEN_2049[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2050 = {1{$random}};
  inputMemBlock_511 = _GEN_2050[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2051 = {1{$random}};
  inputBitsRemaining = _GEN_2051[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2052 = {1{$random}};
  outputMemBlock_0 = _GEN_2052[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2053 = {1{$random}};
  outputMemBlock_1 = _GEN_2053[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2054 = {1{$random}};
  outputMemBlock_2 = _GEN_2054[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2055 = {1{$random}};
  outputMemBlock_3 = _GEN_2055[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2056 = {1{$random}};
  outputMemBlock_4 = _GEN_2056[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2057 = {1{$random}};
  outputMemBlock_5 = _GEN_2057[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2058 = {1{$random}};
  outputMemBlock_6 = _GEN_2058[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2059 = {1{$random}};
  outputMemBlock_7 = _GEN_2059[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2060 = {1{$random}};
  outputMemBlock_8 = _GEN_2060[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2061 = {1{$random}};
  outputMemBlock_9 = _GEN_2061[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2062 = {1{$random}};
  outputMemBlock_10 = _GEN_2062[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2063 = {1{$random}};
  outputMemBlock_11 = _GEN_2063[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2064 = {1{$random}};
  outputMemBlock_12 = _GEN_2064[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2065 = {1{$random}};
  outputMemBlock_13 = _GEN_2065[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2066 = {1{$random}};
  outputMemBlock_14 = _GEN_2066[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2067 = {1{$random}};
  outputMemBlock_15 = _GEN_2067[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2068 = {1{$random}};
  outputMemBlock_16 = _GEN_2068[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2069 = {1{$random}};
  outputMemBlock_17 = _GEN_2069[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2070 = {1{$random}};
  outputMemBlock_18 = _GEN_2070[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2071 = {1{$random}};
  outputMemBlock_19 = _GEN_2071[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2072 = {1{$random}};
  outputMemBlock_20 = _GEN_2072[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2073 = {1{$random}};
  outputMemBlock_21 = _GEN_2073[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2074 = {1{$random}};
  outputMemBlock_22 = _GEN_2074[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2075 = {1{$random}};
  outputMemBlock_23 = _GEN_2075[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2076 = {1{$random}};
  outputMemBlock_24 = _GEN_2076[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2077 = {1{$random}};
  outputMemBlock_25 = _GEN_2077[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2078 = {1{$random}};
  outputMemBlock_26 = _GEN_2078[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2079 = {1{$random}};
  outputMemBlock_27 = _GEN_2079[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2080 = {1{$random}};
  outputMemBlock_28 = _GEN_2080[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2081 = {1{$random}};
  outputMemBlock_29 = _GEN_2081[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2082 = {1{$random}};
  outputMemBlock_30 = _GEN_2082[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2083 = {1{$random}};
  outputMemBlock_31 = _GEN_2083[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2084 = {1{$random}};
  outputMemBlock_32 = _GEN_2084[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2085 = {1{$random}};
  outputMemBlock_33 = _GEN_2085[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2086 = {1{$random}};
  outputMemBlock_34 = _GEN_2086[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2087 = {1{$random}};
  outputMemBlock_35 = _GEN_2087[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2088 = {1{$random}};
  outputMemBlock_36 = _GEN_2088[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2089 = {1{$random}};
  outputMemBlock_37 = _GEN_2089[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2090 = {1{$random}};
  outputMemBlock_38 = _GEN_2090[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2091 = {1{$random}};
  outputMemBlock_39 = _GEN_2091[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2092 = {1{$random}};
  outputMemBlock_40 = _GEN_2092[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2093 = {1{$random}};
  outputMemBlock_41 = _GEN_2093[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2094 = {1{$random}};
  outputMemBlock_42 = _GEN_2094[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2095 = {1{$random}};
  outputMemBlock_43 = _GEN_2095[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2096 = {1{$random}};
  outputMemBlock_44 = _GEN_2096[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2097 = {1{$random}};
  outputMemBlock_45 = _GEN_2097[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2098 = {1{$random}};
  outputMemBlock_46 = _GEN_2098[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2099 = {1{$random}};
  outputMemBlock_47 = _GEN_2099[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2100 = {1{$random}};
  outputMemBlock_48 = _GEN_2100[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2101 = {1{$random}};
  outputMemBlock_49 = _GEN_2101[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2102 = {1{$random}};
  outputMemBlock_50 = _GEN_2102[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2103 = {1{$random}};
  outputMemBlock_51 = _GEN_2103[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2104 = {1{$random}};
  outputMemBlock_52 = _GEN_2104[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2105 = {1{$random}};
  outputMemBlock_53 = _GEN_2105[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2106 = {1{$random}};
  outputMemBlock_54 = _GEN_2106[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2107 = {1{$random}};
  outputMemBlock_55 = _GEN_2107[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2108 = {1{$random}};
  outputMemBlock_56 = _GEN_2108[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2109 = {1{$random}};
  outputMemBlock_57 = _GEN_2109[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2110 = {1{$random}};
  outputMemBlock_58 = _GEN_2110[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2111 = {1{$random}};
  outputMemBlock_59 = _GEN_2111[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2112 = {1{$random}};
  outputMemBlock_60 = _GEN_2112[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2113 = {1{$random}};
  outputMemBlock_61 = _GEN_2113[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2114 = {1{$random}};
  outputMemBlock_62 = _GEN_2114[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2115 = {1{$random}};
  outputMemBlock_63 = _GEN_2115[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2116 = {1{$random}};
  outputMemBlock_64 = _GEN_2116[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2117 = {1{$random}};
  outputMemBlock_65 = _GEN_2117[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2118 = {1{$random}};
  outputMemBlock_66 = _GEN_2118[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2119 = {1{$random}};
  outputMemBlock_67 = _GEN_2119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2120 = {1{$random}};
  outputMemBlock_68 = _GEN_2120[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2121 = {1{$random}};
  outputMemBlock_69 = _GEN_2121[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2122 = {1{$random}};
  outputMemBlock_70 = _GEN_2122[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2123 = {1{$random}};
  outputMemBlock_71 = _GEN_2123[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2124 = {1{$random}};
  outputMemBlock_72 = _GEN_2124[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2125 = {1{$random}};
  outputMemBlock_73 = _GEN_2125[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2126 = {1{$random}};
  outputMemBlock_74 = _GEN_2126[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2127 = {1{$random}};
  outputMemBlock_75 = _GEN_2127[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2128 = {1{$random}};
  outputMemBlock_76 = _GEN_2128[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2129 = {1{$random}};
  outputMemBlock_77 = _GEN_2129[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2130 = {1{$random}};
  outputMemBlock_78 = _GEN_2130[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2131 = {1{$random}};
  outputMemBlock_79 = _GEN_2131[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2132 = {1{$random}};
  outputMemBlock_80 = _GEN_2132[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2133 = {1{$random}};
  outputMemBlock_81 = _GEN_2133[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2134 = {1{$random}};
  outputMemBlock_82 = _GEN_2134[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2135 = {1{$random}};
  outputMemBlock_83 = _GEN_2135[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2136 = {1{$random}};
  outputMemBlock_84 = _GEN_2136[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2137 = {1{$random}};
  outputMemBlock_85 = _GEN_2137[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2138 = {1{$random}};
  outputMemBlock_86 = _GEN_2138[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2139 = {1{$random}};
  outputMemBlock_87 = _GEN_2139[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2140 = {1{$random}};
  outputMemBlock_88 = _GEN_2140[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2141 = {1{$random}};
  outputMemBlock_89 = _GEN_2141[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2142 = {1{$random}};
  outputMemBlock_90 = _GEN_2142[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2143 = {1{$random}};
  outputMemBlock_91 = _GEN_2143[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2144 = {1{$random}};
  outputMemBlock_92 = _GEN_2144[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2145 = {1{$random}};
  outputMemBlock_93 = _GEN_2145[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2146 = {1{$random}};
  outputMemBlock_94 = _GEN_2146[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2147 = {1{$random}};
  outputMemBlock_95 = _GEN_2147[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2148 = {1{$random}};
  outputMemBlock_96 = _GEN_2148[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2149 = {1{$random}};
  outputMemBlock_97 = _GEN_2149[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2150 = {1{$random}};
  outputMemBlock_98 = _GEN_2150[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2151 = {1{$random}};
  outputMemBlock_99 = _GEN_2151[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2152 = {1{$random}};
  outputMemBlock_100 = _GEN_2152[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2153 = {1{$random}};
  outputMemBlock_101 = _GEN_2153[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2154 = {1{$random}};
  outputMemBlock_102 = _GEN_2154[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2155 = {1{$random}};
  outputMemBlock_103 = _GEN_2155[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2156 = {1{$random}};
  outputMemBlock_104 = _GEN_2156[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2157 = {1{$random}};
  outputMemBlock_105 = _GEN_2157[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2158 = {1{$random}};
  outputMemBlock_106 = _GEN_2158[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2159 = {1{$random}};
  outputMemBlock_107 = _GEN_2159[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2160 = {1{$random}};
  outputMemBlock_108 = _GEN_2160[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2161 = {1{$random}};
  outputMemBlock_109 = _GEN_2161[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2162 = {1{$random}};
  outputMemBlock_110 = _GEN_2162[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2163 = {1{$random}};
  outputMemBlock_111 = _GEN_2163[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2164 = {1{$random}};
  outputMemBlock_112 = _GEN_2164[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2165 = {1{$random}};
  outputMemBlock_113 = _GEN_2165[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2166 = {1{$random}};
  outputMemBlock_114 = _GEN_2166[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2167 = {1{$random}};
  outputMemBlock_115 = _GEN_2167[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2168 = {1{$random}};
  outputMemBlock_116 = _GEN_2168[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2169 = {1{$random}};
  outputMemBlock_117 = _GEN_2169[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2170 = {1{$random}};
  outputMemBlock_118 = _GEN_2170[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2171 = {1{$random}};
  outputMemBlock_119 = _GEN_2171[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2172 = {1{$random}};
  outputMemBlock_120 = _GEN_2172[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2173 = {1{$random}};
  outputMemBlock_121 = _GEN_2173[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2174 = {1{$random}};
  outputMemBlock_122 = _GEN_2174[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2175 = {1{$random}};
  outputMemBlock_123 = _GEN_2175[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2176 = {1{$random}};
  outputMemBlock_124 = _GEN_2176[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2177 = {1{$random}};
  outputMemBlock_125 = _GEN_2177[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2178 = {1{$random}};
  outputMemBlock_126 = _GEN_2178[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2179 = {1{$random}};
  outputMemBlock_127 = _GEN_2179[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2180 = {1{$random}};
  outputMemBlock_128 = _GEN_2180[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2181 = {1{$random}};
  outputMemBlock_129 = _GEN_2181[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2182 = {1{$random}};
  outputMemBlock_130 = _GEN_2182[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2183 = {1{$random}};
  outputMemBlock_131 = _GEN_2183[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2184 = {1{$random}};
  outputMemBlock_132 = _GEN_2184[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2185 = {1{$random}};
  outputMemBlock_133 = _GEN_2185[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2186 = {1{$random}};
  outputMemBlock_134 = _GEN_2186[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2187 = {1{$random}};
  outputMemBlock_135 = _GEN_2187[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2188 = {1{$random}};
  outputMemBlock_136 = _GEN_2188[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2189 = {1{$random}};
  outputMemBlock_137 = _GEN_2189[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2190 = {1{$random}};
  outputMemBlock_138 = _GEN_2190[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2191 = {1{$random}};
  outputMemBlock_139 = _GEN_2191[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2192 = {1{$random}};
  outputMemBlock_140 = _GEN_2192[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2193 = {1{$random}};
  outputMemBlock_141 = _GEN_2193[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2194 = {1{$random}};
  outputMemBlock_142 = _GEN_2194[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2195 = {1{$random}};
  outputMemBlock_143 = _GEN_2195[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2196 = {1{$random}};
  outputMemBlock_144 = _GEN_2196[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2197 = {1{$random}};
  outputMemBlock_145 = _GEN_2197[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2198 = {1{$random}};
  outputMemBlock_146 = _GEN_2198[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2199 = {1{$random}};
  outputMemBlock_147 = _GEN_2199[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2200 = {1{$random}};
  outputMemBlock_148 = _GEN_2200[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2201 = {1{$random}};
  outputMemBlock_149 = _GEN_2201[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2202 = {1{$random}};
  outputMemBlock_150 = _GEN_2202[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2203 = {1{$random}};
  outputMemBlock_151 = _GEN_2203[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2204 = {1{$random}};
  outputMemBlock_152 = _GEN_2204[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2205 = {1{$random}};
  outputMemBlock_153 = _GEN_2205[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2206 = {1{$random}};
  outputMemBlock_154 = _GEN_2206[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2207 = {1{$random}};
  outputMemBlock_155 = _GEN_2207[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2208 = {1{$random}};
  outputMemBlock_156 = _GEN_2208[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2209 = {1{$random}};
  outputMemBlock_157 = _GEN_2209[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2210 = {1{$random}};
  outputMemBlock_158 = _GEN_2210[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2211 = {1{$random}};
  outputMemBlock_159 = _GEN_2211[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2212 = {1{$random}};
  outputMemBlock_160 = _GEN_2212[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2213 = {1{$random}};
  outputMemBlock_161 = _GEN_2213[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2214 = {1{$random}};
  outputMemBlock_162 = _GEN_2214[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2215 = {1{$random}};
  outputMemBlock_163 = _GEN_2215[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2216 = {1{$random}};
  outputMemBlock_164 = _GEN_2216[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2217 = {1{$random}};
  outputMemBlock_165 = _GEN_2217[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2218 = {1{$random}};
  outputMemBlock_166 = _GEN_2218[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2219 = {1{$random}};
  outputMemBlock_167 = _GEN_2219[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2220 = {1{$random}};
  outputMemBlock_168 = _GEN_2220[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2221 = {1{$random}};
  outputMemBlock_169 = _GEN_2221[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2222 = {1{$random}};
  outputMemBlock_170 = _GEN_2222[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2223 = {1{$random}};
  outputMemBlock_171 = _GEN_2223[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2224 = {1{$random}};
  outputMemBlock_172 = _GEN_2224[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2225 = {1{$random}};
  outputMemBlock_173 = _GEN_2225[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2226 = {1{$random}};
  outputMemBlock_174 = _GEN_2226[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2227 = {1{$random}};
  outputMemBlock_175 = _GEN_2227[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2228 = {1{$random}};
  outputMemBlock_176 = _GEN_2228[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2229 = {1{$random}};
  outputMemBlock_177 = _GEN_2229[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2230 = {1{$random}};
  outputMemBlock_178 = _GEN_2230[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2231 = {1{$random}};
  outputMemBlock_179 = _GEN_2231[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2232 = {1{$random}};
  outputMemBlock_180 = _GEN_2232[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2233 = {1{$random}};
  outputMemBlock_181 = _GEN_2233[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2234 = {1{$random}};
  outputMemBlock_182 = _GEN_2234[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2235 = {1{$random}};
  outputMemBlock_183 = _GEN_2235[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2236 = {1{$random}};
  outputMemBlock_184 = _GEN_2236[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2237 = {1{$random}};
  outputMemBlock_185 = _GEN_2237[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2238 = {1{$random}};
  outputMemBlock_186 = _GEN_2238[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2239 = {1{$random}};
  outputMemBlock_187 = _GEN_2239[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2240 = {1{$random}};
  outputMemBlock_188 = _GEN_2240[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2241 = {1{$random}};
  outputMemBlock_189 = _GEN_2241[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2242 = {1{$random}};
  outputMemBlock_190 = _GEN_2242[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2243 = {1{$random}};
  outputMemBlock_191 = _GEN_2243[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2244 = {1{$random}};
  outputMemBlock_192 = _GEN_2244[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2245 = {1{$random}};
  outputMemBlock_193 = _GEN_2245[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2246 = {1{$random}};
  outputMemBlock_194 = _GEN_2246[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2247 = {1{$random}};
  outputMemBlock_195 = _GEN_2247[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2248 = {1{$random}};
  outputMemBlock_196 = _GEN_2248[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2249 = {1{$random}};
  outputMemBlock_197 = _GEN_2249[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2250 = {1{$random}};
  outputMemBlock_198 = _GEN_2250[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2251 = {1{$random}};
  outputMemBlock_199 = _GEN_2251[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2252 = {1{$random}};
  outputMemBlock_200 = _GEN_2252[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2253 = {1{$random}};
  outputMemBlock_201 = _GEN_2253[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2254 = {1{$random}};
  outputMemBlock_202 = _GEN_2254[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2255 = {1{$random}};
  outputMemBlock_203 = _GEN_2255[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2256 = {1{$random}};
  outputMemBlock_204 = _GEN_2256[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2257 = {1{$random}};
  outputMemBlock_205 = _GEN_2257[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2258 = {1{$random}};
  outputMemBlock_206 = _GEN_2258[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2259 = {1{$random}};
  outputMemBlock_207 = _GEN_2259[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2260 = {1{$random}};
  outputMemBlock_208 = _GEN_2260[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2261 = {1{$random}};
  outputMemBlock_209 = _GEN_2261[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2262 = {1{$random}};
  outputMemBlock_210 = _GEN_2262[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2263 = {1{$random}};
  outputMemBlock_211 = _GEN_2263[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2264 = {1{$random}};
  outputMemBlock_212 = _GEN_2264[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2265 = {1{$random}};
  outputMemBlock_213 = _GEN_2265[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2266 = {1{$random}};
  outputMemBlock_214 = _GEN_2266[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2267 = {1{$random}};
  outputMemBlock_215 = _GEN_2267[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2268 = {1{$random}};
  outputMemBlock_216 = _GEN_2268[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2269 = {1{$random}};
  outputMemBlock_217 = _GEN_2269[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2270 = {1{$random}};
  outputMemBlock_218 = _GEN_2270[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2271 = {1{$random}};
  outputMemBlock_219 = _GEN_2271[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2272 = {1{$random}};
  outputMemBlock_220 = _GEN_2272[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2273 = {1{$random}};
  outputMemBlock_221 = _GEN_2273[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2274 = {1{$random}};
  outputMemBlock_222 = _GEN_2274[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2275 = {1{$random}};
  outputMemBlock_223 = _GEN_2275[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2276 = {1{$random}};
  outputMemBlock_224 = _GEN_2276[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2277 = {1{$random}};
  outputMemBlock_225 = _GEN_2277[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2278 = {1{$random}};
  outputMemBlock_226 = _GEN_2278[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2279 = {1{$random}};
  outputMemBlock_227 = _GEN_2279[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2280 = {1{$random}};
  outputMemBlock_228 = _GEN_2280[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2281 = {1{$random}};
  outputMemBlock_229 = _GEN_2281[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2282 = {1{$random}};
  outputMemBlock_230 = _GEN_2282[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2283 = {1{$random}};
  outputMemBlock_231 = _GEN_2283[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2284 = {1{$random}};
  outputMemBlock_232 = _GEN_2284[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2285 = {1{$random}};
  outputMemBlock_233 = _GEN_2285[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2286 = {1{$random}};
  outputMemBlock_234 = _GEN_2286[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2287 = {1{$random}};
  outputMemBlock_235 = _GEN_2287[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2288 = {1{$random}};
  outputMemBlock_236 = _GEN_2288[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2289 = {1{$random}};
  outputMemBlock_237 = _GEN_2289[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2290 = {1{$random}};
  outputMemBlock_238 = _GEN_2290[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2291 = {1{$random}};
  outputMemBlock_239 = _GEN_2291[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2292 = {1{$random}};
  outputMemBlock_240 = _GEN_2292[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2293 = {1{$random}};
  outputMemBlock_241 = _GEN_2293[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2294 = {1{$random}};
  outputMemBlock_242 = _GEN_2294[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2295 = {1{$random}};
  outputMemBlock_243 = _GEN_2295[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2296 = {1{$random}};
  outputMemBlock_244 = _GEN_2296[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2297 = {1{$random}};
  outputMemBlock_245 = _GEN_2297[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2298 = {1{$random}};
  outputMemBlock_246 = _GEN_2298[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2299 = {1{$random}};
  outputMemBlock_247 = _GEN_2299[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2300 = {1{$random}};
  outputMemBlock_248 = _GEN_2300[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2301 = {1{$random}};
  outputMemBlock_249 = _GEN_2301[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2302 = {1{$random}};
  outputMemBlock_250 = _GEN_2302[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2303 = {1{$random}};
  outputMemBlock_251 = _GEN_2303[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2304 = {1{$random}};
  outputMemBlock_252 = _GEN_2304[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2305 = {1{$random}};
  outputMemBlock_253 = _GEN_2305[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2306 = {1{$random}};
  outputMemBlock_254 = _GEN_2306[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2307 = {1{$random}};
  outputMemBlock_255 = _GEN_2307[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2308 = {1{$random}};
  outputMemBlock_256 = _GEN_2308[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2309 = {1{$random}};
  outputMemBlock_257 = _GEN_2309[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2310 = {1{$random}};
  outputMemBlock_258 = _GEN_2310[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2311 = {1{$random}};
  outputMemBlock_259 = _GEN_2311[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2312 = {1{$random}};
  outputMemBlock_260 = _GEN_2312[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2313 = {1{$random}};
  outputMemBlock_261 = _GEN_2313[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2314 = {1{$random}};
  outputMemBlock_262 = _GEN_2314[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2315 = {1{$random}};
  outputMemBlock_263 = _GEN_2315[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2316 = {1{$random}};
  outputMemBlock_264 = _GEN_2316[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2317 = {1{$random}};
  outputMemBlock_265 = _GEN_2317[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2318 = {1{$random}};
  outputMemBlock_266 = _GEN_2318[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2319 = {1{$random}};
  outputMemBlock_267 = _GEN_2319[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2320 = {1{$random}};
  outputMemBlock_268 = _GEN_2320[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2321 = {1{$random}};
  outputMemBlock_269 = _GEN_2321[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2322 = {1{$random}};
  outputMemBlock_270 = _GEN_2322[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2323 = {1{$random}};
  outputMemBlock_271 = _GEN_2323[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2324 = {1{$random}};
  outputMemBlock_272 = _GEN_2324[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2325 = {1{$random}};
  outputMemBlock_273 = _GEN_2325[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2326 = {1{$random}};
  outputMemBlock_274 = _GEN_2326[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2327 = {1{$random}};
  outputMemBlock_275 = _GEN_2327[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2328 = {1{$random}};
  outputMemBlock_276 = _GEN_2328[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2329 = {1{$random}};
  outputMemBlock_277 = _GEN_2329[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2330 = {1{$random}};
  outputMemBlock_278 = _GEN_2330[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2331 = {1{$random}};
  outputMemBlock_279 = _GEN_2331[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2332 = {1{$random}};
  outputMemBlock_280 = _GEN_2332[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2333 = {1{$random}};
  outputMemBlock_281 = _GEN_2333[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2334 = {1{$random}};
  outputMemBlock_282 = _GEN_2334[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2335 = {1{$random}};
  outputMemBlock_283 = _GEN_2335[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2336 = {1{$random}};
  outputMemBlock_284 = _GEN_2336[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2337 = {1{$random}};
  outputMemBlock_285 = _GEN_2337[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2338 = {1{$random}};
  outputMemBlock_286 = _GEN_2338[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2339 = {1{$random}};
  outputMemBlock_287 = _GEN_2339[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2340 = {1{$random}};
  outputMemBlock_288 = _GEN_2340[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2341 = {1{$random}};
  outputMemBlock_289 = _GEN_2341[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2342 = {1{$random}};
  outputMemBlock_290 = _GEN_2342[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2343 = {1{$random}};
  outputMemBlock_291 = _GEN_2343[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2344 = {1{$random}};
  outputMemBlock_292 = _GEN_2344[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2345 = {1{$random}};
  outputMemBlock_293 = _GEN_2345[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2346 = {1{$random}};
  outputMemBlock_294 = _GEN_2346[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2347 = {1{$random}};
  outputMemBlock_295 = _GEN_2347[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2348 = {1{$random}};
  outputMemBlock_296 = _GEN_2348[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2349 = {1{$random}};
  outputMemBlock_297 = _GEN_2349[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2350 = {1{$random}};
  outputMemBlock_298 = _GEN_2350[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2351 = {1{$random}};
  outputMemBlock_299 = _GEN_2351[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2352 = {1{$random}};
  outputMemBlock_300 = _GEN_2352[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2353 = {1{$random}};
  outputMemBlock_301 = _GEN_2353[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2354 = {1{$random}};
  outputMemBlock_302 = _GEN_2354[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2355 = {1{$random}};
  outputMemBlock_303 = _GEN_2355[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2356 = {1{$random}};
  outputMemBlock_304 = _GEN_2356[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2357 = {1{$random}};
  outputMemBlock_305 = _GEN_2357[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2358 = {1{$random}};
  outputMemBlock_306 = _GEN_2358[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2359 = {1{$random}};
  outputMemBlock_307 = _GEN_2359[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2360 = {1{$random}};
  outputMemBlock_308 = _GEN_2360[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2361 = {1{$random}};
  outputMemBlock_309 = _GEN_2361[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2362 = {1{$random}};
  outputMemBlock_310 = _GEN_2362[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2363 = {1{$random}};
  outputMemBlock_311 = _GEN_2363[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2364 = {1{$random}};
  outputMemBlock_312 = _GEN_2364[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2365 = {1{$random}};
  outputMemBlock_313 = _GEN_2365[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2366 = {1{$random}};
  outputMemBlock_314 = _GEN_2366[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2367 = {1{$random}};
  outputMemBlock_315 = _GEN_2367[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2368 = {1{$random}};
  outputMemBlock_316 = _GEN_2368[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2369 = {1{$random}};
  outputMemBlock_317 = _GEN_2369[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2370 = {1{$random}};
  outputMemBlock_318 = _GEN_2370[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2371 = {1{$random}};
  outputMemBlock_319 = _GEN_2371[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2372 = {1{$random}};
  outputMemBlock_320 = _GEN_2372[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2373 = {1{$random}};
  outputMemBlock_321 = _GEN_2373[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2374 = {1{$random}};
  outputMemBlock_322 = _GEN_2374[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2375 = {1{$random}};
  outputMemBlock_323 = _GEN_2375[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2376 = {1{$random}};
  outputMemBlock_324 = _GEN_2376[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2377 = {1{$random}};
  outputMemBlock_325 = _GEN_2377[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2378 = {1{$random}};
  outputMemBlock_326 = _GEN_2378[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2379 = {1{$random}};
  outputMemBlock_327 = _GEN_2379[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2380 = {1{$random}};
  outputMemBlock_328 = _GEN_2380[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2381 = {1{$random}};
  outputMemBlock_329 = _GEN_2381[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2382 = {1{$random}};
  outputMemBlock_330 = _GEN_2382[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2383 = {1{$random}};
  outputMemBlock_331 = _GEN_2383[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2384 = {1{$random}};
  outputMemBlock_332 = _GEN_2384[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2385 = {1{$random}};
  outputMemBlock_333 = _GEN_2385[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2386 = {1{$random}};
  outputMemBlock_334 = _GEN_2386[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2387 = {1{$random}};
  outputMemBlock_335 = _GEN_2387[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2388 = {1{$random}};
  outputMemBlock_336 = _GEN_2388[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2389 = {1{$random}};
  outputMemBlock_337 = _GEN_2389[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2390 = {1{$random}};
  outputMemBlock_338 = _GEN_2390[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2391 = {1{$random}};
  outputMemBlock_339 = _GEN_2391[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2392 = {1{$random}};
  outputMemBlock_340 = _GEN_2392[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2393 = {1{$random}};
  outputMemBlock_341 = _GEN_2393[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2394 = {1{$random}};
  outputMemBlock_342 = _GEN_2394[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2395 = {1{$random}};
  outputMemBlock_343 = _GEN_2395[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2396 = {1{$random}};
  outputMemBlock_344 = _GEN_2396[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2397 = {1{$random}};
  outputMemBlock_345 = _GEN_2397[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2398 = {1{$random}};
  outputMemBlock_346 = _GEN_2398[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2399 = {1{$random}};
  outputMemBlock_347 = _GEN_2399[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2400 = {1{$random}};
  outputMemBlock_348 = _GEN_2400[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2401 = {1{$random}};
  outputMemBlock_349 = _GEN_2401[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2402 = {1{$random}};
  outputMemBlock_350 = _GEN_2402[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2403 = {1{$random}};
  outputMemBlock_351 = _GEN_2403[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2404 = {1{$random}};
  outputMemBlock_352 = _GEN_2404[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2405 = {1{$random}};
  outputMemBlock_353 = _GEN_2405[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2406 = {1{$random}};
  outputMemBlock_354 = _GEN_2406[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2407 = {1{$random}};
  outputMemBlock_355 = _GEN_2407[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2408 = {1{$random}};
  outputMemBlock_356 = _GEN_2408[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2409 = {1{$random}};
  outputMemBlock_357 = _GEN_2409[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2410 = {1{$random}};
  outputMemBlock_358 = _GEN_2410[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2411 = {1{$random}};
  outputMemBlock_359 = _GEN_2411[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2412 = {1{$random}};
  outputMemBlock_360 = _GEN_2412[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2413 = {1{$random}};
  outputMemBlock_361 = _GEN_2413[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2414 = {1{$random}};
  outputMemBlock_362 = _GEN_2414[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2415 = {1{$random}};
  outputMemBlock_363 = _GEN_2415[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2416 = {1{$random}};
  outputMemBlock_364 = _GEN_2416[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2417 = {1{$random}};
  outputMemBlock_365 = _GEN_2417[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2418 = {1{$random}};
  outputMemBlock_366 = _GEN_2418[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2419 = {1{$random}};
  outputMemBlock_367 = _GEN_2419[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2420 = {1{$random}};
  outputMemBlock_368 = _GEN_2420[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2421 = {1{$random}};
  outputMemBlock_369 = _GEN_2421[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2422 = {1{$random}};
  outputMemBlock_370 = _GEN_2422[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2423 = {1{$random}};
  outputMemBlock_371 = _GEN_2423[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2424 = {1{$random}};
  outputMemBlock_372 = _GEN_2424[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2425 = {1{$random}};
  outputMemBlock_373 = _GEN_2425[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2426 = {1{$random}};
  outputMemBlock_374 = _GEN_2426[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2427 = {1{$random}};
  outputMemBlock_375 = _GEN_2427[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2428 = {1{$random}};
  outputMemBlock_376 = _GEN_2428[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2429 = {1{$random}};
  outputMemBlock_377 = _GEN_2429[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2430 = {1{$random}};
  outputMemBlock_378 = _GEN_2430[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2431 = {1{$random}};
  outputMemBlock_379 = _GEN_2431[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2432 = {1{$random}};
  outputMemBlock_380 = _GEN_2432[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2433 = {1{$random}};
  outputMemBlock_381 = _GEN_2433[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2434 = {1{$random}};
  outputMemBlock_382 = _GEN_2434[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2435 = {1{$random}};
  outputMemBlock_383 = _GEN_2435[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2436 = {1{$random}};
  outputMemBlock_384 = _GEN_2436[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2437 = {1{$random}};
  outputMemBlock_385 = _GEN_2437[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2438 = {1{$random}};
  outputMemBlock_386 = _GEN_2438[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2439 = {1{$random}};
  outputMemBlock_387 = _GEN_2439[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2440 = {1{$random}};
  outputMemBlock_388 = _GEN_2440[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2441 = {1{$random}};
  outputMemBlock_389 = _GEN_2441[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2442 = {1{$random}};
  outputMemBlock_390 = _GEN_2442[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2443 = {1{$random}};
  outputMemBlock_391 = _GEN_2443[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2444 = {1{$random}};
  outputMemBlock_392 = _GEN_2444[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2445 = {1{$random}};
  outputMemBlock_393 = _GEN_2445[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2446 = {1{$random}};
  outputMemBlock_394 = _GEN_2446[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2447 = {1{$random}};
  outputMemBlock_395 = _GEN_2447[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2448 = {1{$random}};
  outputMemBlock_396 = _GEN_2448[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2449 = {1{$random}};
  outputMemBlock_397 = _GEN_2449[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2450 = {1{$random}};
  outputMemBlock_398 = _GEN_2450[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2451 = {1{$random}};
  outputMemBlock_399 = _GEN_2451[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2452 = {1{$random}};
  outputMemBlock_400 = _GEN_2452[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2453 = {1{$random}};
  outputMemBlock_401 = _GEN_2453[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2454 = {1{$random}};
  outputMemBlock_402 = _GEN_2454[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2455 = {1{$random}};
  outputMemBlock_403 = _GEN_2455[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2456 = {1{$random}};
  outputMemBlock_404 = _GEN_2456[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2457 = {1{$random}};
  outputMemBlock_405 = _GEN_2457[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2458 = {1{$random}};
  outputMemBlock_406 = _GEN_2458[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2459 = {1{$random}};
  outputMemBlock_407 = _GEN_2459[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2460 = {1{$random}};
  outputMemBlock_408 = _GEN_2460[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2461 = {1{$random}};
  outputMemBlock_409 = _GEN_2461[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2462 = {1{$random}};
  outputMemBlock_410 = _GEN_2462[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2463 = {1{$random}};
  outputMemBlock_411 = _GEN_2463[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2464 = {1{$random}};
  outputMemBlock_412 = _GEN_2464[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2465 = {1{$random}};
  outputMemBlock_413 = _GEN_2465[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2466 = {1{$random}};
  outputMemBlock_414 = _GEN_2466[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2467 = {1{$random}};
  outputMemBlock_415 = _GEN_2467[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2468 = {1{$random}};
  outputMemBlock_416 = _GEN_2468[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2469 = {1{$random}};
  outputMemBlock_417 = _GEN_2469[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2470 = {1{$random}};
  outputMemBlock_418 = _GEN_2470[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2471 = {1{$random}};
  outputMemBlock_419 = _GEN_2471[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2472 = {1{$random}};
  outputMemBlock_420 = _GEN_2472[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2473 = {1{$random}};
  outputMemBlock_421 = _GEN_2473[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2474 = {1{$random}};
  outputMemBlock_422 = _GEN_2474[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2475 = {1{$random}};
  outputMemBlock_423 = _GEN_2475[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2476 = {1{$random}};
  outputMemBlock_424 = _GEN_2476[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2477 = {1{$random}};
  outputMemBlock_425 = _GEN_2477[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2478 = {1{$random}};
  outputMemBlock_426 = _GEN_2478[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2479 = {1{$random}};
  outputMemBlock_427 = _GEN_2479[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2480 = {1{$random}};
  outputMemBlock_428 = _GEN_2480[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2481 = {1{$random}};
  outputMemBlock_429 = _GEN_2481[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2482 = {1{$random}};
  outputMemBlock_430 = _GEN_2482[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2483 = {1{$random}};
  outputMemBlock_431 = _GEN_2483[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2484 = {1{$random}};
  outputMemBlock_432 = _GEN_2484[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2485 = {1{$random}};
  outputMemBlock_433 = _GEN_2485[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2486 = {1{$random}};
  outputMemBlock_434 = _GEN_2486[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2487 = {1{$random}};
  outputMemBlock_435 = _GEN_2487[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2488 = {1{$random}};
  outputMemBlock_436 = _GEN_2488[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2489 = {1{$random}};
  outputMemBlock_437 = _GEN_2489[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2490 = {1{$random}};
  outputMemBlock_438 = _GEN_2490[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2491 = {1{$random}};
  outputMemBlock_439 = _GEN_2491[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2492 = {1{$random}};
  outputMemBlock_440 = _GEN_2492[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2493 = {1{$random}};
  outputMemBlock_441 = _GEN_2493[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2494 = {1{$random}};
  outputMemBlock_442 = _GEN_2494[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2495 = {1{$random}};
  outputMemBlock_443 = _GEN_2495[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2496 = {1{$random}};
  outputMemBlock_444 = _GEN_2496[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2497 = {1{$random}};
  outputMemBlock_445 = _GEN_2497[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2498 = {1{$random}};
  outputMemBlock_446 = _GEN_2498[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2499 = {1{$random}};
  outputMemBlock_447 = _GEN_2499[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2500 = {1{$random}};
  outputMemBlock_448 = _GEN_2500[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2501 = {1{$random}};
  outputMemBlock_449 = _GEN_2501[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2502 = {1{$random}};
  outputMemBlock_450 = _GEN_2502[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2503 = {1{$random}};
  outputMemBlock_451 = _GEN_2503[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2504 = {1{$random}};
  outputMemBlock_452 = _GEN_2504[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2505 = {1{$random}};
  outputMemBlock_453 = _GEN_2505[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2506 = {1{$random}};
  outputMemBlock_454 = _GEN_2506[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2507 = {1{$random}};
  outputMemBlock_455 = _GEN_2507[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2508 = {1{$random}};
  outputMemBlock_456 = _GEN_2508[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2509 = {1{$random}};
  outputMemBlock_457 = _GEN_2509[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2510 = {1{$random}};
  outputMemBlock_458 = _GEN_2510[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2511 = {1{$random}};
  outputMemBlock_459 = _GEN_2511[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2512 = {1{$random}};
  outputMemBlock_460 = _GEN_2512[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2513 = {1{$random}};
  outputMemBlock_461 = _GEN_2513[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2514 = {1{$random}};
  outputMemBlock_462 = _GEN_2514[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2515 = {1{$random}};
  outputMemBlock_463 = _GEN_2515[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2516 = {1{$random}};
  outputMemBlock_464 = _GEN_2516[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2517 = {1{$random}};
  outputMemBlock_465 = _GEN_2517[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2518 = {1{$random}};
  outputMemBlock_466 = _GEN_2518[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2519 = {1{$random}};
  outputMemBlock_467 = _GEN_2519[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2520 = {1{$random}};
  outputMemBlock_468 = _GEN_2520[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2521 = {1{$random}};
  outputMemBlock_469 = _GEN_2521[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2522 = {1{$random}};
  outputMemBlock_470 = _GEN_2522[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2523 = {1{$random}};
  outputMemBlock_471 = _GEN_2523[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2524 = {1{$random}};
  outputMemBlock_472 = _GEN_2524[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2525 = {1{$random}};
  outputMemBlock_473 = _GEN_2525[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2526 = {1{$random}};
  outputMemBlock_474 = _GEN_2526[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2527 = {1{$random}};
  outputMemBlock_475 = _GEN_2527[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2528 = {1{$random}};
  outputMemBlock_476 = _GEN_2528[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2529 = {1{$random}};
  outputMemBlock_477 = _GEN_2529[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2530 = {1{$random}};
  outputMemBlock_478 = _GEN_2530[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2531 = {1{$random}};
  outputMemBlock_479 = _GEN_2531[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2532 = {1{$random}};
  outputMemBlock_480 = _GEN_2532[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2533 = {1{$random}};
  outputMemBlock_481 = _GEN_2533[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2534 = {1{$random}};
  outputMemBlock_482 = _GEN_2534[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2535 = {1{$random}};
  outputMemBlock_483 = _GEN_2535[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2536 = {1{$random}};
  outputMemBlock_484 = _GEN_2536[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2537 = {1{$random}};
  outputMemBlock_485 = _GEN_2537[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2538 = {1{$random}};
  outputMemBlock_486 = _GEN_2538[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2539 = {1{$random}};
  outputMemBlock_487 = _GEN_2539[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2540 = {1{$random}};
  outputMemBlock_488 = _GEN_2540[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2541 = {1{$random}};
  outputMemBlock_489 = _GEN_2541[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2542 = {1{$random}};
  outputMemBlock_490 = _GEN_2542[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2543 = {1{$random}};
  outputMemBlock_491 = _GEN_2543[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2544 = {1{$random}};
  outputMemBlock_492 = _GEN_2544[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2545 = {1{$random}};
  outputMemBlock_493 = _GEN_2545[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2546 = {1{$random}};
  outputMemBlock_494 = _GEN_2546[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2547 = {1{$random}};
  outputMemBlock_495 = _GEN_2547[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2548 = {1{$random}};
  outputMemBlock_496 = _GEN_2548[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2549 = {1{$random}};
  outputMemBlock_497 = _GEN_2549[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2550 = {1{$random}};
  outputMemBlock_498 = _GEN_2550[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2551 = {1{$random}};
  outputMemBlock_499 = _GEN_2551[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2552 = {1{$random}};
  outputMemBlock_500 = _GEN_2552[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2553 = {1{$random}};
  outputMemBlock_501 = _GEN_2553[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2554 = {1{$random}};
  outputMemBlock_502 = _GEN_2554[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2555 = {1{$random}};
  outputMemBlock_503 = _GEN_2555[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2556 = {1{$random}};
  outputMemBlock_504 = _GEN_2556[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2557 = {1{$random}};
  outputMemBlock_505 = _GEN_2557[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2558 = {1{$random}};
  outputMemBlock_506 = _GEN_2558[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2559 = {1{$random}};
  outputMemBlock_507 = _GEN_2559[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2560 = {1{$random}};
  outputMemBlock_508 = _GEN_2560[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2561 = {1{$random}};
  outputMemBlock_509 = _GEN_2561[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2562 = {1{$random}};
  outputMemBlock_510 = _GEN_2562[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2563 = {1{$random}};
  outputMemBlock_511 = _GEN_2563[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2564 = {1{$random}};
  outputBits = _GEN_2564[9:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (inputAdvance) begin
      inputMemBlock_0 <= inputMemBlock_1;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_0 <= _T_540;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_1 <= inputMemBlock_2;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_1 <= _T_541;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_2 <= inputMemBlock_3;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_2 <= _T_542;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_3 <= inputMemBlock_4;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_3 <= _T_543;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_4 <= inputMemBlock_5;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_4 <= _T_544;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_5 <= inputMemBlock_6;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_5 <= _T_545;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_6 <= inputMemBlock_7;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_6 <= _T_546;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_7 <= inputMemBlock_8;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_7 <= _T_547;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_8 <= inputMemBlock_9;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_8 <= _T_548;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_9 <= inputMemBlock_10;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_9 <= _T_549;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_10 <= inputMemBlock_11;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_10 <= _T_550;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_11 <= inputMemBlock_12;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_11 <= _T_551;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_12 <= inputMemBlock_13;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_12 <= _T_552;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_13 <= inputMemBlock_14;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_13 <= _T_553;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_14 <= inputMemBlock_15;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_14 <= _T_554;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_15 <= inputMemBlock_16;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_15 <= _T_555;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_16 <= inputMemBlock_17;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_16 <= _T_556;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_17 <= inputMemBlock_18;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_17 <= _T_557;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_18 <= inputMemBlock_19;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_18 <= _T_558;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_19 <= inputMemBlock_20;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_19 <= _T_559;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_20 <= inputMemBlock_21;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_20 <= _T_560;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_21 <= inputMemBlock_22;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_21 <= _T_561;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_22 <= inputMemBlock_23;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_22 <= _T_562;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_23 <= inputMemBlock_24;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_23 <= _T_563;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_24 <= inputMemBlock_25;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_24 <= _T_564;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_25 <= inputMemBlock_26;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_25 <= _T_565;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_26 <= inputMemBlock_27;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_26 <= _T_566;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_27 <= inputMemBlock_28;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_27 <= _T_567;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_28 <= inputMemBlock_29;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_28 <= _T_568;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_29 <= inputMemBlock_30;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_29 <= _T_569;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_30 <= inputMemBlock_31;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_30 <= _T_570;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_31 <= inputMemBlock_32;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_31 <= _T_571;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_32 <= inputMemBlock_33;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_32 <= _T_572;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_33 <= inputMemBlock_34;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_33 <= _T_573;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_34 <= inputMemBlock_35;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_34 <= _T_574;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_35 <= inputMemBlock_36;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_35 <= _T_575;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_36 <= inputMemBlock_37;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_36 <= _T_576;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_37 <= inputMemBlock_38;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_37 <= _T_577;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_38 <= inputMemBlock_39;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_38 <= _T_578;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_39 <= inputMemBlock_40;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_39 <= _T_579;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_40 <= inputMemBlock_41;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_40 <= _T_580;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_41 <= inputMemBlock_42;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_41 <= _T_581;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_42 <= inputMemBlock_43;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_42 <= _T_582;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_43 <= inputMemBlock_44;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_43 <= _T_583;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_44 <= inputMemBlock_45;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_44 <= _T_584;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_45 <= inputMemBlock_46;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_45 <= _T_585;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_46 <= inputMemBlock_47;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_46 <= _T_586;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_47 <= inputMemBlock_48;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_47 <= _T_587;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_48 <= inputMemBlock_49;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_48 <= _T_588;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_49 <= inputMemBlock_50;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_49 <= _T_589;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_50 <= inputMemBlock_51;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_50 <= _T_590;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_51 <= inputMemBlock_52;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_51 <= _T_591;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_52 <= inputMemBlock_53;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_52 <= _T_592;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_53 <= inputMemBlock_54;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_53 <= _T_593;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_54 <= inputMemBlock_55;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_54 <= _T_594;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_55 <= inputMemBlock_56;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_55 <= _T_595;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_56 <= inputMemBlock_57;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_56 <= _T_596;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_57 <= inputMemBlock_58;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_57 <= _T_597;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_58 <= inputMemBlock_59;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_58 <= _T_598;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_59 <= inputMemBlock_60;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_59 <= _T_599;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_60 <= inputMemBlock_61;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_60 <= _T_600;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_61 <= inputMemBlock_62;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_61 <= _T_601;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_62 <= inputMemBlock_63;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_62 <= _T_602;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_63 <= inputMemBlock_64;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_63 <= _T_603;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_64 <= inputMemBlock_65;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_64 <= _T_604;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_65 <= inputMemBlock_66;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_65 <= _T_605;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_66 <= inputMemBlock_67;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_66 <= _T_606;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_67 <= inputMemBlock_68;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_67 <= _T_607;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_68 <= inputMemBlock_69;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_68 <= _T_608;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_69 <= inputMemBlock_70;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_69 <= _T_609;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_70 <= inputMemBlock_71;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_70 <= _T_610;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_71 <= inputMemBlock_72;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_71 <= _T_611;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_72 <= inputMemBlock_73;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_72 <= _T_612;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_73 <= inputMemBlock_74;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_73 <= _T_613;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_74 <= inputMemBlock_75;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_74 <= _T_614;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_75 <= inputMemBlock_76;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_75 <= _T_615;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_76 <= inputMemBlock_77;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_76 <= _T_616;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_77 <= inputMemBlock_78;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_77 <= _T_617;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_78 <= inputMemBlock_79;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_78 <= _T_618;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_79 <= inputMemBlock_80;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_79 <= _T_619;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_80 <= inputMemBlock_81;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_80 <= _T_620;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_81 <= inputMemBlock_82;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_81 <= _T_621;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_82 <= inputMemBlock_83;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_82 <= _T_622;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_83 <= inputMemBlock_84;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_83 <= _T_623;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_84 <= inputMemBlock_85;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_84 <= _T_624;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_85 <= inputMemBlock_86;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_85 <= _T_625;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_86 <= inputMemBlock_87;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_86 <= _T_626;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_87 <= inputMemBlock_88;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_87 <= _T_627;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_88 <= inputMemBlock_89;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_88 <= _T_628;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_89 <= inputMemBlock_90;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_89 <= _T_629;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_90 <= inputMemBlock_91;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_90 <= _T_630;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_91 <= inputMemBlock_92;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_91 <= _T_631;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_92 <= inputMemBlock_93;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_92 <= _T_632;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_93 <= inputMemBlock_94;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_93 <= _T_633;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_94 <= inputMemBlock_95;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_94 <= _T_634;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_95 <= inputMemBlock_96;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_95 <= _T_635;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_96 <= inputMemBlock_97;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_96 <= _T_636;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_97 <= inputMemBlock_98;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_97 <= _T_637;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_98 <= inputMemBlock_99;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_98 <= _T_638;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_99 <= inputMemBlock_100;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_99 <= _T_639;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_100 <= inputMemBlock_101;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_100 <= _T_640;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_101 <= inputMemBlock_102;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_101 <= _T_641;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_102 <= inputMemBlock_103;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_102 <= _T_642;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_103 <= inputMemBlock_104;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_103 <= _T_643;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_104 <= inputMemBlock_105;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_104 <= _T_644;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_105 <= inputMemBlock_106;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_105 <= _T_645;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_106 <= inputMemBlock_107;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_106 <= _T_646;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_107 <= inputMemBlock_108;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_107 <= _T_647;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_108 <= inputMemBlock_109;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_108 <= _T_648;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_109 <= inputMemBlock_110;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_109 <= _T_649;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_110 <= inputMemBlock_111;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_110 <= _T_650;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_111 <= inputMemBlock_112;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_111 <= _T_651;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_112 <= inputMemBlock_113;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_112 <= _T_652;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_113 <= inputMemBlock_114;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_113 <= _T_653;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_114 <= inputMemBlock_115;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_114 <= _T_654;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_115 <= inputMemBlock_116;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_115 <= _T_655;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_116 <= inputMemBlock_117;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_116 <= _T_656;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_117 <= inputMemBlock_118;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_117 <= _T_657;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_118 <= inputMemBlock_119;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_118 <= _T_658;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_119 <= inputMemBlock_120;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_119 <= _T_659;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_120 <= inputMemBlock_121;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_120 <= _T_660;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_121 <= inputMemBlock_122;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_121 <= _T_661;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_122 <= inputMemBlock_123;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_122 <= _T_662;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_123 <= inputMemBlock_124;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_123 <= _T_663;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_124 <= inputMemBlock_125;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_124 <= _T_664;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_125 <= inputMemBlock_126;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_125 <= _T_665;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_126 <= inputMemBlock_127;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_126 <= _T_666;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_127 <= inputMemBlock_128;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_127 <= _T_667;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_128 <= inputMemBlock_129;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_128 <= _T_668;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_129 <= inputMemBlock_130;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_129 <= _T_669;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_130 <= inputMemBlock_131;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_130 <= _T_670;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_131 <= inputMemBlock_132;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_131 <= _T_671;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_132 <= inputMemBlock_133;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_132 <= _T_672;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_133 <= inputMemBlock_134;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_133 <= _T_673;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_134 <= inputMemBlock_135;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_134 <= _T_674;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_135 <= inputMemBlock_136;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_135 <= _T_675;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_136 <= inputMemBlock_137;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_136 <= _T_676;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_137 <= inputMemBlock_138;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_137 <= _T_677;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_138 <= inputMemBlock_139;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_138 <= _T_678;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_139 <= inputMemBlock_140;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_139 <= _T_679;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_140 <= inputMemBlock_141;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_140 <= _T_680;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_141 <= inputMemBlock_142;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_141 <= _T_681;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_142 <= inputMemBlock_143;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_142 <= _T_682;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_143 <= inputMemBlock_144;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_143 <= _T_683;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_144 <= inputMemBlock_145;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_144 <= _T_684;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_145 <= inputMemBlock_146;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_145 <= _T_685;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_146 <= inputMemBlock_147;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_146 <= _T_686;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_147 <= inputMemBlock_148;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_147 <= _T_687;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_148 <= inputMemBlock_149;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_148 <= _T_688;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_149 <= inputMemBlock_150;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_149 <= _T_689;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_150 <= inputMemBlock_151;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_150 <= _T_690;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_151 <= inputMemBlock_152;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_151 <= _T_691;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_152 <= inputMemBlock_153;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_152 <= _T_692;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_153 <= inputMemBlock_154;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_153 <= _T_693;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_154 <= inputMemBlock_155;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_154 <= _T_694;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_155 <= inputMemBlock_156;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_155 <= _T_695;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_156 <= inputMemBlock_157;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_156 <= _T_696;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_157 <= inputMemBlock_158;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_157 <= _T_697;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_158 <= inputMemBlock_159;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_158 <= _T_698;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_159 <= inputMemBlock_160;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_159 <= _T_699;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_160 <= inputMemBlock_161;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_160 <= _T_700;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_161 <= inputMemBlock_162;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_161 <= _T_701;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_162 <= inputMemBlock_163;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_162 <= _T_702;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_163 <= inputMemBlock_164;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_163 <= _T_703;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_164 <= inputMemBlock_165;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_164 <= _T_704;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_165 <= inputMemBlock_166;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_165 <= _T_705;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_166 <= inputMemBlock_167;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_166 <= _T_706;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_167 <= inputMemBlock_168;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_167 <= _T_707;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_168 <= inputMemBlock_169;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_168 <= _T_708;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_169 <= inputMemBlock_170;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_169 <= _T_709;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_170 <= inputMemBlock_171;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_170 <= _T_710;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_171 <= inputMemBlock_172;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_171 <= _T_711;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_172 <= inputMemBlock_173;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_172 <= _T_712;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_173 <= inputMemBlock_174;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_173 <= _T_713;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_174 <= inputMemBlock_175;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_174 <= _T_714;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_175 <= inputMemBlock_176;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_175 <= _T_715;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_176 <= inputMemBlock_177;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_176 <= _T_716;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_177 <= inputMemBlock_178;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_177 <= _T_717;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_178 <= inputMemBlock_179;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_178 <= _T_718;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_179 <= inputMemBlock_180;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_179 <= _T_719;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_180 <= inputMemBlock_181;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_180 <= _T_720;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_181 <= inputMemBlock_182;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_181 <= _T_721;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_182 <= inputMemBlock_183;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_182 <= _T_722;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_183 <= inputMemBlock_184;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_183 <= _T_723;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_184 <= inputMemBlock_185;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_184 <= _T_724;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_185 <= inputMemBlock_186;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_185 <= _T_725;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_186 <= inputMemBlock_187;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_186 <= _T_726;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_187 <= inputMemBlock_188;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_187 <= _T_727;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_188 <= inputMemBlock_189;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_188 <= _T_728;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_189 <= inputMemBlock_190;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_189 <= _T_729;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_190 <= inputMemBlock_191;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_190 <= _T_730;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_191 <= inputMemBlock_192;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_191 <= _T_731;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_192 <= inputMemBlock_193;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_192 <= _T_732;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_193 <= inputMemBlock_194;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_193 <= _T_733;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_194 <= inputMemBlock_195;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_194 <= _T_734;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_195 <= inputMemBlock_196;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_195 <= _T_735;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_196 <= inputMemBlock_197;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_196 <= _T_736;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_197 <= inputMemBlock_198;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_197 <= _T_737;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_198 <= inputMemBlock_199;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_198 <= _T_738;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_199 <= inputMemBlock_200;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_199 <= _T_739;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_200 <= inputMemBlock_201;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_200 <= _T_740;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_201 <= inputMemBlock_202;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_201 <= _T_741;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_202 <= inputMemBlock_203;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_202 <= _T_742;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_203 <= inputMemBlock_204;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_203 <= _T_743;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_204 <= inputMemBlock_205;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_204 <= _T_744;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_205 <= inputMemBlock_206;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_205 <= _T_745;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_206 <= inputMemBlock_207;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_206 <= _T_746;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_207 <= inputMemBlock_208;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_207 <= _T_747;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_208 <= inputMemBlock_209;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_208 <= _T_748;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_209 <= inputMemBlock_210;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_209 <= _T_749;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_210 <= inputMemBlock_211;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_210 <= _T_750;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_211 <= inputMemBlock_212;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_211 <= _T_751;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_212 <= inputMemBlock_213;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_212 <= _T_752;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_213 <= inputMemBlock_214;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_213 <= _T_753;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_214 <= inputMemBlock_215;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_214 <= _T_754;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_215 <= inputMemBlock_216;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_215 <= _T_755;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_216 <= inputMemBlock_217;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_216 <= _T_756;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_217 <= inputMemBlock_218;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_217 <= _T_757;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_218 <= inputMemBlock_219;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_218 <= _T_758;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_219 <= inputMemBlock_220;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_219 <= _T_759;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_220 <= inputMemBlock_221;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_220 <= _T_760;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_221 <= inputMemBlock_222;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_221 <= _T_761;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_222 <= inputMemBlock_223;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_222 <= _T_762;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_223 <= inputMemBlock_224;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_223 <= _T_763;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_224 <= inputMemBlock_225;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_224 <= _T_764;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_225 <= inputMemBlock_226;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_225 <= _T_765;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_226 <= inputMemBlock_227;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_226 <= _T_766;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_227 <= inputMemBlock_228;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_227 <= _T_767;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_228 <= inputMemBlock_229;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_228 <= _T_768;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_229 <= inputMemBlock_230;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_229 <= _T_769;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_230 <= inputMemBlock_231;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_230 <= _T_770;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_231 <= inputMemBlock_232;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_231 <= _T_771;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_232 <= inputMemBlock_233;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_232 <= _T_772;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_233 <= inputMemBlock_234;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_233 <= _T_773;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_234 <= inputMemBlock_235;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_234 <= _T_774;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_235 <= inputMemBlock_236;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_235 <= _T_775;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_236 <= inputMemBlock_237;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_236 <= _T_776;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_237 <= inputMemBlock_238;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_237 <= _T_777;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_238 <= inputMemBlock_239;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_238 <= _T_778;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_239 <= inputMemBlock_240;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_239 <= _T_779;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_240 <= inputMemBlock_241;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_240 <= _T_780;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_241 <= inputMemBlock_242;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_241 <= _T_781;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_242 <= inputMemBlock_243;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_242 <= _T_782;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_243 <= inputMemBlock_244;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_243 <= _T_783;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_244 <= inputMemBlock_245;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_244 <= _T_784;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_245 <= inputMemBlock_246;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_245 <= _T_785;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_246 <= inputMemBlock_247;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_246 <= _T_786;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_247 <= inputMemBlock_248;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_247 <= _T_787;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_248 <= inputMemBlock_249;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_248 <= _T_788;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_249 <= inputMemBlock_250;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_249 <= _T_789;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_250 <= inputMemBlock_251;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_250 <= _T_790;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_251 <= inputMemBlock_252;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_251 <= _T_791;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_252 <= inputMemBlock_253;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_252 <= _T_792;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_253 <= inputMemBlock_254;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_253 <= _T_793;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_254 <= inputMemBlock_255;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_254 <= _T_794;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_255 <= inputMemBlock_256;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_255 <= _T_795;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_256 <= inputMemBlock_257;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_256 <= _T_796;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_257 <= inputMemBlock_258;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_257 <= _T_797;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_258 <= inputMemBlock_259;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_258 <= _T_798;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_259 <= inputMemBlock_260;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_259 <= _T_799;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_260 <= inputMemBlock_261;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_260 <= _T_800;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_261 <= inputMemBlock_262;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_261 <= _T_801;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_262 <= inputMemBlock_263;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_262 <= _T_802;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_263 <= inputMemBlock_264;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_263 <= _T_803;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_264 <= inputMemBlock_265;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_264 <= _T_804;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_265 <= inputMemBlock_266;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_265 <= _T_805;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_266 <= inputMemBlock_267;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_266 <= _T_806;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_267 <= inputMemBlock_268;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_267 <= _T_807;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_268 <= inputMemBlock_269;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_268 <= _T_808;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_269 <= inputMemBlock_270;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_269 <= _T_809;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_270 <= inputMemBlock_271;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_270 <= _T_810;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_271 <= inputMemBlock_272;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_271 <= _T_811;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_272 <= inputMemBlock_273;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_272 <= _T_812;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_273 <= inputMemBlock_274;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_273 <= _T_813;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_274 <= inputMemBlock_275;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_274 <= _T_814;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_275 <= inputMemBlock_276;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_275 <= _T_815;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_276 <= inputMemBlock_277;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_276 <= _T_816;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_277 <= inputMemBlock_278;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_277 <= _T_817;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_278 <= inputMemBlock_279;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_278 <= _T_818;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_279 <= inputMemBlock_280;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_279 <= _T_819;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_280 <= inputMemBlock_281;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_280 <= _T_820;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_281 <= inputMemBlock_282;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_281 <= _T_821;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_282 <= inputMemBlock_283;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_282 <= _T_822;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_283 <= inputMemBlock_284;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_283 <= _T_823;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_284 <= inputMemBlock_285;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_284 <= _T_824;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_285 <= inputMemBlock_286;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_285 <= _T_825;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_286 <= inputMemBlock_287;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_286 <= _T_826;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_287 <= inputMemBlock_288;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_287 <= _T_827;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_288 <= inputMemBlock_289;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_288 <= _T_828;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_289 <= inputMemBlock_290;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_289 <= _T_829;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_290 <= inputMemBlock_291;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_290 <= _T_830;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_291 <= inputMemBlock_292;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_291 <= _T_831;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_292 <= inputMemBlock_293;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_292 <= _T_832;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_293 <= inputMemBlock_294;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_293 <= _T_833;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_294 <= inputMemBlock_295;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_294 <= _T_834;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_295 <= inputMemBlock_296;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_295 <= _T_835;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_296 <= inputMemBlock_297;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_296 <= _T_836;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_297 <= inputMemBlock_298;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_297 <= _T_837;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_298 <= inputMemBlock_299;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_298 <= _T_838;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_299 <= inputMemBlock_300;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_299 <= _T_839;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_300 <= inputMemBlock_301;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_300 <= _T_840;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_301 <= inputMemBlock_302;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_301 <= _T_841;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_302 <= inputMemBlock_303;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_302 <= _T_842;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_303 <= inputMemBlock_304;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_303 <= _T_843;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_304 <= inputMemBlock_305;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_304 <= _T_844;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_305 <= inputMemBlock_306;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_305 <= _T_845;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_306 <= inputMemBlock_307;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_306 <= _T_846;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_307 <= inputMemBlock_308;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_307 <= _T_847;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_308 <= inputMemBlock_309;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_308 <= _T_848;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_309 <= inputMemBlock_310;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_309 <= _T_849;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_310 <= inputMemBlock_311;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_310 <= _T_850;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_311 <= inputMemBlock_312;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_311 <= _T_851;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_312 <= inputMemBlock_313;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_312 <= _T_852;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_313 <= inputMemBlock_314;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_313 <= _T_853;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_314 <= inputMemBlock_315;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_314 <= _T_854;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_315 <= inputMemBlock_316;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_315 <= _T_855;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_316 <= inputMemBlock_317;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_316 <= _T_856;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_317 <= inputMemBlock_318;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_317 <= _T_857;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_318 <= inputMemBlock_319;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_318 <= _T_858;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_319 <= inputMemBlock_320;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_319 <= _T_859;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_320 <= inputMemBlock_321;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_320 <= _T_860;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_321 <= inputMemBlock_322;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_321 <= _T_861;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_322 <= inputMemBlock_323;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_322 <= _T_862;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_323 <= inputMemBlock_324;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_323 <= _T_863;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_324 <= inputMemBlock_325;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_324 <= _T_864;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_325 <= inputMemBlock_326;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_325 <= _T_865;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_326 <= inputMemBlock_327;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_326 <= _T_866;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_327 <= inputMemBlock_328;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_327 <= _T_867;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_328 <= inputMemBlock_329;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_328 <= _T_868;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_329 <= inputMemBlock_330;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_329 <= _T_869;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_330 <= inputMemBlock_331;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_330 <= _T_870;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_331 <= inputMemBlock_332;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_331 <= _T_871;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_332 <= inputMemBlock_333;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_332 <= _T_872;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_333 <= inputMemBlock_334;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_333 <= _T_873;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_334 <= inputMemBlock_335;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_334 <= _T_874;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_335 <= inputMemBlock_336;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_335 <= _T_875;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_336 <= inputMemBlock_337;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_336 <= _T_876;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_337 <= inputMemBlock_338;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_337 <= _T_877;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_338 <= inputMemBlock_339;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_338 <= _T_878;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_339 <= inputMemBlock_340;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_339 <= _T_879;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_340 <= inputMemBlock_341;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_340 <= _T_880;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_341 <= inputMemBlock_342;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_341 <= _T_881;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_342 <= inputMemBlock_343;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_342 <= _T_882;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_343 <= inputMemBlock_344;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_343 <= _T_883;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_344 <= inputMemBlock_345;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_344 <= _T_884;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_345 <= inputMemBlock_346;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_345 <= _T_885;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_346 <= inputMemBlock_347;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_346 <= _T_886;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_347 <= inputMemBlock_348;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_347 <= _T_887;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_348 <= inputMemBlock_349;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_348 <= _T_888;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_349 <= inputMemBlock_350;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_349 <= _T_889;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_350 <= inputMemBlock_351;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_350 <= _T_890;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_351 <= inputMemBlock_352;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_351 <= _T_891;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_352 <= inputMemBlock_353;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_352 <= _T_892;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_353 <= inputMemBlock_354;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_353 <= _T_893;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_354 <= inputMemBlock_355;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_354 <= _T_894;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_355 <= inputMemBlock_356;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_355 <= _T_895;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_356 <= inputMemBlock_357;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_356 <= _T_896;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_357 <= inputMemBlock_358;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_357 <= _T_897;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_358 <= inputMemBlock_359;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_358 <= _T_898;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_359 <= inputMemBlock_360;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_359 <= _T_899;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_360 <= inputMemBlock_361;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_360 <= _T_900;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_361 <= inputMemBlock_362;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_361 <= _T_901;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_362 <= inputMemBlock_363;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_362 <= _T_902;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_363 <= inputMemBlock_364;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_363 <= _T_903;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_364 <= inputMemBlock_365;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_364 <= _T_904;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_365 <= inputMemBlock_366;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_365 <= _T_905;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_366 <= inputMemBlock_367;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_366 <= _T_906;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_367 <= inputMemBlock_368;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_367 <= _T_907;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_368 <= inputMemBlock_369;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_368 <= _T_908;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_369 <= inputMemBlock_370;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_369 <= _T_909;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_370 <= inputMemBlock_371;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_370 <= _T_910;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_371 <= inputMemBlock_372;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_371 <= _T_911;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_372 <= inputMemBlock_373;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_372 <= _T_912;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_373 <= inputMemBlock_374;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_373 <= _T_913;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_374 <= inputMemBlock_375;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_374 <= _T_914;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_375 <= inputMemBlock_376;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_375 <= _T_915;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_376 <= inputMemBlock_377;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_376 <= _T_916;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_377 <= inputMemBlock_378;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_377 <= _T_917;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_378 <= inputMemBlock_379;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_378 <= _T_918;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_379 <= inputMemBlock_380;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_379 <= _T_919;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_380 <= inputMemBlock_381;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_380 <= _T_920;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_381 <= inputMemBlock_382;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_381 <= _T_921;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_382 <= inputMemBlock_383;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_382 <= _T_922;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_383 <= inputMemBlock_384;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_383 <= _T_923;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_384 <= inputMemBlock_385;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_384 <= _T_924;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_385 <= inputMemBlock_386;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_385 <= _T_925;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_386 <= inputMemBlock_387;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_386 <= _T_926;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_387 <= inputMemBlock_388;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_387 <= _T_927;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_388 <= inputMemBlock_389;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_388 <= _T_928;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_389 <= inputMemBlock_390;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_389 <= _T_929;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_390 <= inputMemBlock_391;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_390 <= _T_930;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_391 <= inputMemBlock_392;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_391 <= _T_931;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_392 <= inputMemBlock_393;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_392 <= _T_932;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_393 <= inputMemBlock_394;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_393 <= _T_933;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_394 <= inputMemBlock_395;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_394 <= _T_934;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_395 <= inputMemBlock_396;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_395 <= _T_935;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_396 <= inputMemBlock_397;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_396 <= _T_936;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_397 <= inputMemBlock_398;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_397 <= _T_937;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_398 <= inputMemBlock_399;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_398 <= _T_938;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_399 <= inputMemBlock_400;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_399 <= _T_939;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_400 <= inputMemBlock_401;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_400 <= _T_940;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_401 <= inputMemBlock_402;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_401 <= _T_941;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_402 <= inputMemBlock_403;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_402 <= _T_942;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_403 <= inputMemBlock_404;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_403 <= _T_943;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_404 <= inputMemBlock_405;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_404 <= _T_944;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_405 <= inputMemBlock_406;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_405 <= _T_945;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_406 <= inputMemBlock_407;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_406 <= _T_946;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_407 <= inputMemBlock_408;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_407 <= _T_947;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_408 <= inputMemBlock_409;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_408 <= _T_948;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_409 <= inputMemBlock_410;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_409 <= _T_949;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_410 <= inputMemBlock_411;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_410 <= _T_950;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_411 <= inputMemBlock_412;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_411 <= _T_951;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_412 <= inputMemBlock_413;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_412 <= _T_952;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_413 <= inputMemBlock_414;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_413 <= _T_953;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_414 <= inputMemBlock_415;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_414 <= _T_954;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_415 <= inputMemBlock_416;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_415 <= _T_955;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_416 <= inputMemBlock_417;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_416 <= _T_956;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_417 <= inputMemBlock_418;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_417 <= _T_957;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_418 <= inputMemBlock_419;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_418 <= _T_958;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_419 <= inputMemBlock_420;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_419 <= _T_959;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_420 <= inputMemBlock_421;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_420 <= _T_960;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_421 <= inputMemBlock_422;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_421 <= _T_961;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_422 <= inputMemBlock_423;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_422 <= _T_962;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_423 <= inputMemBlock_424;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_423 <= _T_963;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_424 <= inputMemBlock_425;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_424 <= _T_964;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_425 <= inputMemBlock_426;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_425 <= _T_965;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_426 <= inputMemBlock_427;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_426 <= _T_966;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_427 <= inputMemBlock_428;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_427 <= _T_967;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_428 <= inputMemBlock_429;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_428 <= _T_968;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_429 <= inputMemBlock_430;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_429 <= _T_969;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_430 <= inputMemBlock_431;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_430 <= _T_970;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_431 <= inputMemBlock_432;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_431 <= _T_971;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_432 <= inputMemBlock_433;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_432 <= _T_972;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_433 <= inputMemBlock_434;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_433 <= _T_973;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_434 <= inputMemBlock_435;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_434 <= _T_974;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_435 <= inputMemBlock_436;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_435 <= _T_975;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_436 <= inputMemBlock_437;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_436 <= _T_976;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_437 <= inputMemBlock_438;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_437 <= _T_977;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_438 <= inputMemBlock_439;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_438 <= _T_978;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_439 <= inputMemBlock_440;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_439 <= _T_979;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_440 <= inputMemBlock_441;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_440 <= _T_980;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_441 <= inputMemBlock_442;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_441 <= _T_981;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_442 <= inputMemBlock_443;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_442 <= _T_982;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_443 <= inputMemBlock_444;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_443 <= _T_983;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_444 <= inputMemBlock_445;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_444 <= _T_984;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_445 <= inputMemBlock_446;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_445 <= _T_985;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_446 <= inputMemBlock_447;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_446 <= _T_986;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_447 <= inputMemBlock_448;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_447 <= _T_987;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_448 <= inputMemBlock_449;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_448 <= _T_988;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_449 <= inputMemBlock_450;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_449 <= _T_989;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_450 <= inputMemBlock_451;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_450 <= _T_990;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_451 <= inputMemBlock_452;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_451 <= _T_991;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_452 <= inputMemBlock_453;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_452 <= _T_992;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_453 <= inputMemBlock_454;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_453 <= _T_993;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_454 <= inputMemBlock_455;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_454 <= _T_994;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_455 <= inputMemBlock_456;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_455 <= _T_995;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_456 <= inputMemBlock_457;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_456 <= _T_996;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_457 <= inputMemBlock_458;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_457 <= _T_997;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_458 <= inputMemBlock_459;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_458 <= _T_998;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_459 <= inputMemBlock_460;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_459 <= _T_999;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_460 <= inputMemBlock_461;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_460 <= _T_1000;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_461 <= inputMemBlock_462;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_461 <= _T_1001;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_462 <= inputMemBlock_463;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_462 <= _T_1002;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_463 <= inputMemBlock_464;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_463 <= _T_1003;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_464 <= inputMemBlock_465;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_464 <= _T_1004;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_465 <= inputMemBlock_466;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_465 <= _T_1005;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_466 <= inputMemBlock_467;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_466 <= _T_1006;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_467 <= inputMemBlock_468;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_467 <= _T_1007;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_468 <= inputMemBlock_469;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_468 <= _T_1008;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_469 <= inputMemBlock_470;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_469 <= _T_1009;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_470 <= inputMemBlock_471;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_470 <= _T_1010;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_471 <= inputMemBlock_472;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_471 <= _T_1011;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_472 <= inputMemBlock_473;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_472 <= _T_1012;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_473 <= inputMemBlock_474;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_473 <= _T_1013;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_474 <= inputMemBlock_475;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_474 <= _T_1014;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_475 <= inputMemBlock_476;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_475 <= _T_1015;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_476 <= inputMemBlock_477;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_476 <= _T_1016;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_477 <= inputMemBlock_478;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_477 <= _T_1017;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_478 <= inputMemBlock_479;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_478 <= _T_1018;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_479 <= inputMemBlock_480;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_479 <= _T_1019;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_480 <= inputMemBlock_481;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_480 <= _T_1020;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_481 <= inputMemBlock_482;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_481 <= _T_1021;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_482 <= inputMemBlock_483;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_482 <= _T_1022;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_483 <= inputMemBlock_484;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_483 <= _T_1023;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_484 <= inputMemBlock_485;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_484 <= _T_1024;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_485 <= inputMemBlock_486;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_485 <= _T_1025;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_486 <= inputMemBlock_487;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_486 <= _T_1026;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_487 <= inputMemBlock_488;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_487 <= _T_1027;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_488 <= inputMemBlock_489;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_488 <= _T_1028;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_489 <= inputMemBlock_490;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_489 <= _T_1029;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_490 <= inputMemBlock_491;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_490 <= _T_1030;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_491 <= inputMemBlock_492;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_491 <= _T_1031;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_492 <= inputMemBlock_493;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_492 <= _T_1032;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_493 <= inputMemBlock_494;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_493 <= _T_1033;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_494 <= inputMemBlock_495;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_494 <= _T_1034;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_495 <= inputMemBlock_496;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_495 <= _T_1035;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_496 <= inputMemBlock_497;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_496 <= _T_1036;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_497 <= inputMemBlock_498;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_497 <= _T_1037;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_498 <= inputMemBlock_499;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_498 <= _T_1038;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_499 <= inputMemBlock_500;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_499 <= _T_1039;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_500 <= inputMemBlock_501;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_500 <= _T_1040;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_501 <= inputMemBlock_502;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_501 <= _T_1041;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_502 <= inputMemBlock_503;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_502 <= _T_1042;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_503 <= inputMemBlock_504;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_503 <= _T_1043;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_504 <= inputMemBlock_505;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_504 <= _T_1044;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_505 <= inputMemBlock_506;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_505 <= _T_1045;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_506 <= inputMemBlock_507;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_506 <= _T_1046;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_507 <= inputMemBlock_508;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_507 <= _T_1047;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_508 <= inputMemBlock_509;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_508 <= _T_1048;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_509 <= inputMemBlock_510;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_509 <= _T_1049;
      end
    end
    if (inputAdvance) begin
      inputMemBlock_510 <= inputMemBlock_511;
    end else begin
      if (io_inputMemBlockValid) begin
        inputMemBlock_510 <= _T_1050;
      end
    end
    if (io_inputMemBlockValid) begin
      inputMemBlock_511 <= _T_1051;
    end
    if (reset) begin
      inputBitsRemaining <= 10'h0;
    end else begin
      if (inputAdvance) begin
        inputBitsRemaining <= _T_1585;
      end else begin
        if (io_inputMemBlockValid) begin
          inputBitsRemaining <= io_inputBits;
        end
      end
    end
    if (nextBitValid) begin
      outputMemBlock_0 <= outputMemBlock_1;
    end
    if (nextBitValid) begin
      outputMemBlock_1 <= outputMemBlock_2;
    end
    if (nextBitValid) begin
      outputMemBlock_2 <= outputMemBlock_3;
    end
    if (nextBitValid) begin
      outputMemBlock_3 <= outputMemBlock_4;
    end
    if (nextBitValid) begin
      outputMemBlock_4 <= outputMemBlock_5;
    end
    if (nextBitValid) begin
      outputMemBlock_5 <= outputMemBlock_6;
    end
    if (nextBitValid) begin
      outputMemBlock_6 <= outputMemBlock_7;
    end
    if (nextBitValid) begin
      outputMemBlock_7 <= outputMemBlock_8;
    end
    if (nextBitValid) begin
      outputMemBlock_8 <= outputMemBlock_9;
    end
    if (nextBitValid) begin
      outputMemBlock_9 <= outputMemBlock_10;
    end
    if (nextBitValid) begin
      outputMemBlock_10 <= outputMemBlock_11;
    end
    if (nextBitValid) begin
      outputMemBlock_11 <= outputMemBlock_12;
    end
    if (nextBitValid) begin
      outputMemBlock_12 <= outputMemBlock_13;
    end
    if (nextBitValid) begin
      outputMemBlock_13 <= outputMemBlock_14;
    end
    if (nextBitValid) begin
      outputMemBlock_14 <= outputMemBlock_15;
    end
    if (nextBitValid) begin
      outputMemBlock_15 <= outputMemBlock_16;
    end
    if (nextBitValid) begin
      outputMemBlock_16 <= outputMemBlock_17;
    end
    if (nextBitValid) begin
      outputMemBlock_17 <= outputMemBlock_18;
    end
    if (nextBitValid) begin
      outputMemBlock_18 <= outputMemBlock_19;
    end
    if (nextBitValid) begin
      outputMemBlock_19 <= outputMemBlock_20;
    end
    if (nextBitValid) begin
      outputMemBlock_20 <= outputMemBlock_21;
    end
    if (nextBitValid) begin
      outputMemBlock_21 <= outputMemBlock_22;
    end
    if (nextBitValid) begin
      outputMemBlock_22 <= outputMemBlock_23;
    end
    if (nextBitValid) begin
      outputMemBlock_23 <= outputMemBlock_24;
    end
    if (nextBitValid) begin
      outputMemBlock_24 <= outputMemBlock_25;
    end
    if (nextBitValid) begin
      outputMemBlock_25 <= outputMemBlock_26;
    end
    if (nextBitValid) begin
      outputMemBlock_26 <= outputMemBlock_27;
    end
    if (nextBitValid) begin
      outputMemBlock_27 <= outputMemBlock_28;
    end
    if (nextBitValid) begin
      outputMemBlock_28 <= outputMemBlock_29;
    end
    if (nextBitValid) begin
      outputMemBlock_29 <= outputMemBlock_30;
    end
    if (nextBitValid) begin
      outputMemBlock_30 <= outputMemBlock_31;
    end
    if (nextBitValid) begin
      outputMemBlock_31 <= outputMemBlock_32;
    end
    if (nextBitValid) begin
      outputMemBlock_32 <= outputMemBlock_33;
    end
    if (nextBitValid) begin
      outputMemBlock_33 <= outputMemBlock_34;
    end
    if (nextBitValid) begin
      outputMemBlock_34 <= outputMemBlock_35;
    end
    if (nextBitValid) begin
      outputMemBlock_35 <= outputMemBlock_36;
    end
    if (nextBitValid) begin
      outputMemBlock_36 <= outputMemBlock_37;
    end
    if (nextBitValid) begin
      outputMemBlock_37 <= outputMemBlock_38;
    end
    if (nextBitValid) begin
      outputMemBlock_38 <= outputMemBlock_39;
    end
    if (nextBitValid) begin
      outputMemBlock_39 <= outputMemBlock_40;
    end
    if (nextBitValid) begin
      outputMemBlock_40 <= outputMemBlock_41;
    end
    if (nextBitValid) begin
      outputMemBlock_41 <= outputMemBlock_42;
    end
    if (nextBitValid) begin
      outputMemBlock_42 <= outputMemBlock_43;
    end
    if (nextBitValid) begin
      outputMemBlock_43 <= outputMemBlock_44;
    end
    if (nextBitValid) begin
      outputMemBlock_44 <= outputMemBlock_45;
    end
    if (nextBitValid) begin
      outputMemBlock_45 <= outputMemBlock_46;
    end
    if (nextBitValid) begin
      outputMemBlock_46 <= outputMemBlock_47;
    end
    if (nextBitValid) begin
      outputMemBlock_47 <= outputMemBlock_48;
    end
    if (nextBitValid) begin
      outputMemBlock_48 <= outputMemBlock_49;
    end
    if (nextBitValid) begin
      outputMemBlock_49 <= outputMemBlock_50;
    end
    if (nextBitValid) begin
      outputMemBlock_50 <= outputMemBlock_51;
    end
    if (nextBitValid) begin
      outputMemBlock_51 <= outputMemBlock_52;
    end
    if (nextBitValid) begin
      outputMemBlock_52 <= outputMemBlock_53;
    end
    if (nextBitValid) begin
      outputMemBlock_53 <= outputMemBlock_54;
    end
    if (nextBitValid) begin
      outputMemBlock_54 <= outputMemBlock_55;
    end
    if (nextBitValid) begin
      outputMemBlock_55 <= outputMemBlock_56;
    end
    if (nextBitValid) begin
      outputMemBlock_56 <= outputMemBlock_57;
    end
    if (nextBitValid) begin
      outputMemBlock_57 <= outputMemBlock_58;
    end
    if (nextBitValid) begin
      outputMemBlock_58 <= outputMemBlock_59;
    end
    if (nextBitValid) begin
      outputMemBlock_59 <= outputMemBlock_60;
    end
    if (nextBitValid) begin
      outputMemBlock_60 <= outputMemBlock_61;
    end
    if (nextBitValid) begin
      outputMemBlock_61 <= outputMemBlock_62;
    end
    if (nextBitValid) begin
      outputMemBlock_62 <= outputMemBlock_63;
    end
    if (nextBitValid) begin
      outputMemBlock_63 <= outputMemBlock_64;
    end
    if (nextBitValid) begin
      outputMemBlock_64 <= outputMemBlock_65;
    end
    if (nextBitValid) begin
      outputMemBlock_65 <= outputMemBlock_66;
    end
    if (nextBitValid) begin
      outputMemBlock_66 <= outputMemBlock_67;
    end
    if (nextBitValid) begin
      outputMemBlock_67 <= outputMemBlock_68;
    end
    if (nextBitValid) begin
      outputMemBlock_68 <= outputMemBlock_69;
    end
    if (nextBitValid) begin
      outputMemBlock_69 <= outputMemBlock_70;
    end
    if (nextBitValid) begin
      outputMemBlock_70 <= outputMemBlock_71;
    end
    if (nextBitValid) begin
      outputMemBlock_71 <= outputMemBlock_72;
    end
    if (nextBitValid) begin
      outputMemBlock_72 <= outputMemBlock_73;
    end
    if (nextBitValid) begin
      outputMemBlock_73 <= outputMemBlock_74;
    end
    if (nextBitValid) begin
      outputMemBlock_74 <= outputMemBlock_75;
    end
    if (nextBitValid) begin
      outputMemBlock_75 <= outputMemBlock_76;
    end
    if (nextBitValid) begin
      outputMemBlock_76 <= outputMemBlock_77;
    end
    if (nextBitValid) begin
      outputMemBlock_77 <= outputMemBlock_78;
    end
    if (nextBitValid) begin
      outputMemBlock_78 <= outputMemBlock_79;
    end
    if (nextBitValid) begin
      outputMemBlock_79 <= outputMemBlock_80;
    end
    if (nextBitValid) begin
      outputMemBlock_80 <= outputMemBlock_81;
    end
    if (nextBitValid) begin
      outputMemBlock_81 <= outputMemBlock_82;
    end
    if (nextBitValid) begin
      outputMemBlock_82 <= outputMemBlock_83;
    end
    if (nextBitValid) begin
      outputMemBlock_83 <= outputMemBlock_84;
    end
    if (nextBitValid) begin
      outputMemBlock_84 <= outputMemBlock_85;
    end
    if (nextBitValid) begin
      outputMemBlock_85 <= outputMemBlock_86;
    end
    if (nextBitValid) begin
      outputMemBlock_86 <= outputMemBlock_87;
    end
    if (nextBitValid) begin
      outputMemBlock_87 <= outputMemBlock_88;
    end
    if (nextBitValid) begin
      outputMemBlock_88 <= outputMemBlock_89;
    end
    if (nextBitValid) begin
      outputMemBlock_89 <= outputMemBlock_90;
    end
    if (nextBitValid) begin
      outputMemBlock_90 <= outputMemBlock_91;
    end
    if (nextBitValid) begin
      outputMemBlock_91 <= outputMemBlock_92;
    end
    if (nextBitValid) begin
      outputMemBlock_92 <= outputMemBlock_93;
    end
    if (nextBitValid) begin
      outputMemBlock_93 <= outputMemBlock_94;
    end
    if (nextBitValid) begin
      outputMemBlock_94 <= outputMemBlock_95;
    end
    if (nextBitValid) begin
      outputMemBlock_95 <= outputMemBlock_96;
    end
    if (nextBitValid) begin
      outputMemBlock_96 <= outputMemBlock_97;
    end
    if (nextBitValid) begin
      outputMemBlock_97 <= outputMemBlock_98;
    end
    if (nextBitValid) begin
      outputMemBlock_98 <= outputMemBlock_99;
    end
    if (nextBitValid) begin
      outputMemBlock_99 <= outputMemBlock_100;
    end
    if (nextBitValid) begin
      outputMemBlock_100 <= outputMemBlock_101;
    end
    if (nextBitValid) begin
      outputMemBlock_101 <= outputMemBlock_102;
    end
    if (nextBitValid) begin
      outputMemBlock_102 <= outputMemBlock_103;
    end
    if (nextBitValid) begin
      outputMemBlock_103 <= outputMemBlock_104;
    end
    if (nextBitValid) begin
      outputMemBlock_104 <= outputMemBlock_105;
    end
    if (nextBitValid) begin
      outputMemBlock_105 <= outputMemBlock_106;
    end
    if (nextBitValid) begin
      outputMemBlock_106 <= outputMemBlock_107;
    end
    if (nextBitValid) begin
      outputMemBlock_107 <= outputMemBlock_108;
    end
    if (nextBitValid) begin
      outputMemBlock_108 <= outputMemBlock_109;
    end
    if (nextBitValid) begin
      outputMemBlock_109 <= outputMemBlock_110;
    end
    if (nextBitValid) begin
      outputMemBlock_110 <= outputMemBlock_111;
    end
    if (nextBitValid) begin
      outputMemBlock_111 <= outputMemBlock_112;
    end
    if (nextBitValid) begin
      outputMemBlock_112 <= outputMemBlock_113;
    end
    if (nextBitValid) begin
      outputMemBlock_113 <= outputMemBlock_114;
    end
    if (nextBitValid) begin
      outputMemBlock_114 <= outputMemBlock_115;
    end
    if (nextBitValid) begin
      outputMemBlock_115 <= outputMemBlock_116;
    end
    if (nextBitValid) begin
      outputMemBlock_116 <= outputMemBlock_117;
    end
    if (nextBitValid) begin
      outputMemBlock_117 <= outputMemBlock_118;
    end
    if (nextBitValid) begin
      outputMemBlock_118 <= outputMemBlock_119;
    end
    if (nextBitValid) begin
      outputMemBlock_119 <= outputMemBlock_120;
    end
    if (nextBitValid) begin
      outputMemBlock_120 <= outputMemBlock_121;
    end
    if (nextBitValid) begin
      outputMemBlock_121 <= outputMemBlock_122;
    end
    if (nextBitValid) begin
      outputMemBlock_122 <= outputMemBlock_123;
    end
    if (nextBitValid) begin
      outputMemBlock_123 <= outputMemBlock_124;
    end
    if (nextBitValid) begin
      outputMemBlock_124 <= outputMemBlock_125;
    end
    if (nextBitValid) begin
      outputMemBlock_125 <= outputMemBlock_126;
    end
    if (nextBitValid) begin
      outputMemBlock_126 <= outputMemBlock_127;
    end
    if (nextBitValid) begin
      outputMemBlock_127 <= outputMemBlock_128;
    end
    if (nextBitValid) begin
      outputMemBlock_128 <= outputMemBlock_129;
    end
    if (nextBitValid) begin
      outputMemBlock_129 <= outputMemBlock_130;
    end
    if (nextBitValid) begin
      outputMemBlock_130 <= outputMemBlock_131;
    end
    if (nextBitValid) begin
      outputMemBlock_131 <= outputMemBlock_132;
    end
    if (nextBitValid) begin
      outputMemBlock_132 <= outputMemBlock_133;
    end
    if (nextBitValid) begin
      outputMemBlock_133 <= outputMemBlock_134;
    end
    if (nextBitValid) begin
      outputMemBlock_134 <= outputMemBlock_135;
    end
    if (nextBitValid) begin
      outputMemBlock_135 <= outputMemBlock_136;
    end
    if (nextBitValid) begin
      outputMemBlock_136 <= outputMemBlock_137;
    end
    if (nextBitValid) begin
      outputMemBlock_137 <= outputMemBlock_138;
    end
    if (nextBitValid) begin
      outputMemBlock_138 <= outputMemBlock_139;
    end
    if (nextBitValid) begin
      outputMemBlock_139 <= outputMemBlock_140;
    end
    if (nextBitValid) begin
      outputMemBlock_140 <= outputMemBlock_141;
    end
    if (nextBitValid) begin
      outputMemBlock_141 <= outputMemBlock_142;
    end
    if (nextBitValid) begin
      outputMemBlock_142 <= outputMemBlock_143;
    end
    if (nextBitValid) begin
      outputMemBlock_143 <= outputMemBlock_144;
    end
    if (nextBitValid) begin
      outputMemBlock_144 <= outputMemBlock_145;
    end
    if (nextBitValid) begin
      outputMemBlock_145 <= outputMemBlock_146;
    end
    if (nextBitValid) begin
      outputMemBlock_146 <= outputMemBlock_147;
    end
    if (nextBitValid) begin
      outputMemBlock_147 <= outputMemBlock_148;
    end
    if (nextBitValid) begin
      outputMemBlock_148 <= outputMemBlock_149;
    end
    if (nextBitValid) begin
      outputMemBlock_149 <= outputMemBlock_150;
    end
    if (nextBitValid) begin
      outputMemBlock_150 <= outputMemBlock_151;
    end
    if (nextBitValid) begin
      outputMemBlock_151 <= outputMemBlock_152;
    end
    if (nextBitValid) begin
      outputMemBlock_152 <= outputMemBlock_153;
    end
    if (nextBitValid) begin
      outputMemBlock_153 <= outputMemBlock_154;
    end
    if (nextBitValid) begin
      outputMemBlock_154 <= outputMemBlock_155;
    end
    if (nextBitValid) begin
      outputMemBlock_155 <= outputMemBlock_156;
    end
    if (nextBitValid) begin
      outputMemBlock_156 <= outputMemBlock_157;
    end
    if (nextBitValid) begin
      outputMemBlock_157 <= outputMemBlock_158;
    end
    if (nextBitValid) begin
      outputMemBlock_158 <= outputMemBlock_159;
    end
    if (nextBitValid) begin
      outputMemBlock_159 <= outputMemBlock_160;
    end
    if (nextBitValid) begin
      outputMemBlock_160 <= outputMemBlock_161;
    end
    if (nextBitValid) begin
      outputMemBlock_161 <= outputMemBlock_162;
    end
    if (nextBitValid) begin
      outputMemBlock_162 <= outputMemBlock_163;
    end
    if (nextBitValid) begin
      outputMemBlock_163 <= outputMemBlock_164;
    end
    if (nextBitValid) begin
      outputMemBlock_164 <= outputMemBlock_165;
    end
    if (nextBitValid) begin
      outputMemBlock_165 <= outputMemBlock_166;
    end
    if (nextBitValid) begin
      outputMemBlock_166 <= outputMemBlock_167;
    end
    if (nextBitValid) begin
      outputMemBlock_167 <= outputMemBlock_168;
    end
    if (nextBitValid) begin
      outputMemBlock_168 <= outputMemBlock_169;
    end
    if (nextBitValid) begin
      outputMemBlock_169 <= outputMemBlock_170;
    end
    if (nextBitValid) begin
      outputMemBlock_170 <= outputMemBlock_171;
    end
    if (nextBitValid) begin
      outputMemBlock_171 <= outputMemBlock_172;
    end
    if (nextBitValid) begin
      outputMemBlock_172 <= outputMemBlock_173;
    end
    if (nextBitValid) begin
      outputMemBlock_173 <= outputMemBlock_174;
    end
    if (nextBitValid) begin
      outputMemBlock_174 <= outputMemBlock_175;
    end
    if (nextBitValid) begin
      outputMemBlock_175 <= outputMemBlock_176;
    end
    if (nextBitValid) begin
      outputMemBlock_176 <= outputMemBlock_177;
    end
    if (nextBitValid) begin
      outputMemBlock_177 <= outputMemBlock_178;
    end
    if (nextBitValid) begin
      outputMemBlock_178 <= outputMemBlock_179;
    end
    if (nextBitValid) begin
      outputMemBlock_179 <= outputMemBlock_180;
    end
    if (nextBitValid) begin
      outputMemBlock_180 <= outputMemBlock_181;
    end
    if (nextBitValid) begin
      outputMemBlock_181 <= outputMemBlock_182;
    end
    if (nextBitValid) begin
      outputMemBlock_182 <= outputMemBlock_183;
    end
    if (nextBitValid) begin
      outputMemBlock_183 <= outputMemBlock_184;
    end
    if (nextBitValid) begin
      outputMemBlock_184 <= outputMemBlock_185;
    end
    if (nextBitValid) begin
      outputMemBlock_185 <= outputMemBlock_186;
    end
    if (nextBitValid) begin
      outputMemBlock_186 <= outputMemBlock_187;
    end
    if (nextBitValid) begin
      outputMemBlock_187 <= outputMemBlock_188;
    end
    if (nextBitValid) begin
      outputMemBlock_188 <= outputMemBlock_189;
    end
    if (nextBitValid) begin
      outputMemBlock_189 <= outputMemBlock_190;
    end
    if (nextBitValid) begin
      outputMemBlock_190 <= outputMemBlock_191;
    end
    if (nextBitValid) begin
      outputMemBlock_191 <= outputMemBlock_192;
    end
    if (nextBitValid) begin
      outputMemBlock_192 <= outputMemBlock_193;
    end
    if (nextBitValid) begin
      outputMemBlock_193 <= outputMemBlock_194;
    end
    if (nextBitValid) begin
      outputMemBlock_194 <= outputMemBlock_195;
    end
    if (nextBitValid) begin
      outputMemBlock_195 <= outputMemBlock_196;
    end
    if (nextBitValid) begin
      outputMemBlock_196 <= outputMemBlock_197;
    end
    if (nextBitValid) begin
      outputMemBlock_197 <= outputMemBlock_198;
    end
    if (nextBitValid) begin
      outputMemBlock_198 <= outputMemBlock_199;
    end
    if (nextBitValid) begin
      outputMemBlock_199 <= outputMemBlock_200;
    end
    if (nextBitValid) begin
      outputMemBlock_200 <= outputMemBlock_201;
    end
    if (nextBitValid) begin
      outputMemBlock_201 <= outputMemBlock_202;
    end
    if (nextBitValid) begin
      outputMemBlock_202 <= outputMemBlock_203;
    end
    if (nextBitValid) begin
      outputMemBlock_203 <= outputMemBlock_204;
    end
    if (nextBitValid) begin
      outputMemBlock_204 <= outputMemBlock_205;
    end
    if (nextBitValid) begin
      outputMemBlock_205 <= outputMemBlock_206;
    end
    if (nextBitValid) begin
      outputMemBlock_206 <= outputMemBlock_207;
    end
    if (nextBitValid) begin
      outputMemBlock_207 <= outputMemBlock_208;
    end
    if (nextBitValid) begin
      outputMemBlock_208 <= outputMemBlock_209;
    end
    if (nextBitValid) begin
      outputMemBlock_209 <= outputMemBlock_210;
    end
    if (nextBitValid) begin
      outputMemBlock_210 <= outputMemBlock_211;
    end
    if (nextBitValid) begin
      outputMemBlock_211 <= outputMemBlock_212;
    end
    if (nextBitValid) begin
      outputMemBlock_212 <= outputMemBlock_213;
    end
    if (nextBitValid) begin
      outputMemBlock_213 <= outputMemBlock_214;
    end
    if (nextBitValid) begin
      outputMemBlock_214 <= outputMemBlock_215;
    end
    if (nextBitValid) begin
      outputMemBlock_215 <= outputMemBlock_216;
    end
    if (nextBitValid) begin
      outputMemBlock_216 <= outputMemBlock_217;
    end
    if (nextBitValid) begin
      outputMemBlock_217 <= outputMemBlock_218;
    end
    if (nextBitValid) begin
      outputMemBlock_218 <= outputMemBlock_219;
    end
    if (nextBitValid) begin
      outputMemBlock_219 <= outputMemBlock_220;
    end
    if (nextBitValid) begin
      outputMemBlock_220 <= outputMemBlock_221;
    end
    if (nextBitValid) begin
      outputMemBlock_221 <= outputMemBlock_222;
    end
    if (nextBitValid) begin
      outputMemBlock_222 <= outputMemBlock_223;
    end
    if (nextBitValid) begin
      outputMemBlock_223 <= outputMemBlock_224;
    end
    if (nextBitValid) begin
      outputMemBlock_224 <= outputMemBlock_225;
    end
    if (nextBitValid) begin
      outputMemBlock_225 <= outputMemBlock_226;
    end
    if (nextBitValid) begin
      outputMemBlock_226 <= outputMemBlock_227;
    end
    if (nextBitValid) begin
      outputMemBlock_227 <= outputMemBlock_228;
    end
    if (nextBitValid) begin
      outputMemBlock_228 <= outputMemBlock_229;
    end
    if (nextBitValid) begin
      outputMemBlock_229 <= outputMemBlock_230;
    end
    if (nextBitValid) begin
      outputMemBlock_230 <= outputMemBlock_231;
    end
    if (nextBitValid) begin
      outputMemBlock_231 <= outputMemBlock_232;
    end
    if (nextBitValid) begin
      outputMemBlock_232 <= outputMemBlock_233;
    end
    if (nextBitValid) begin
      outputMemBlock_233 <= outputMemBlock_234;
    end
    if (nextBitValid) begin
      outputMemBlock_234 <= outputMemBlock_235;
    end
    if (nextBitValid) begin
      outputMemBlock_235 <= outputMemBlock_236;
    end
    if (nextBitValid) begin
      outputMemBlock_236 <= outputMemBlock_237;
    end
    if (nextBitValid) begin
      outputMemBlock_237 <= outputMemBlock_238;
    end
    if (nextBitValid) begin
      outputMemBlock_238 <= outputMemBlock_239;
    end
    if (nextBitValid) begin
      outputMemBlock_239 <= outputMemBlock_240;
    end
    if (nextBitValid) begin
      outputMemBlock_240 <= outputMemBlock_241;
    end
    if (nextBitValid) begin
      outputMemBlock_241 <= outputMemBlock_242;
    end
    if (nextBitValid) begin
      outputMemBlock_242 <= outputMemBlock_243;
    end
    if (nextBitValid) begin
      outputMemBlock_243 <= outputMemBlock_244;
    end
    if (nextBitValid) begin
      outputMemBlock_244 <= outputMemBlock_245;
    end
    if (nextBitValid) begin
      outputMemBlock_245 <= outputMemBlock_246;
    end
    if (nextBitValid) begin
      outputMemBlock_246 <= outputMemBlock_247;
    end
    if (nextBitValid) begin
      outputMemBlock_247 <= outputMemBlock_248;
    end
    if (nextBitValid) begin
      outputMemBlock_248 <= outputMemBlock_249;
    end
    if (nextBitValid) begin
      outputMemBlock_249 <= outputMemBlock_250;
    end
    if (nextBitValid) begin
      outputMemBlock_250 <= outputMemBlock_251;
    end
    if (nextBitValid) begin
      outputMemBlock_251 <= outputMemBlock_252;
    end
    if (nextBitValid) begin
      outputMemBlock_252 <= outputMemBlock_253;
    end
    if (nextBitValid) begin
      outputMemBlock_253 <= outputMemBlock_254;
    end
    if (nextBitValid) begin
      outputMemBlock_254 <= outputMemBlock_255;
    end
    if (nextBitValid) begin
      outputMemBlock_255 <= outputMemBlock_256;
    end
    if (nextBitValid) begin
      outputMemBlock_256 <= outputMemBlock_257;
    end
    if (nextBitValid) begin
      outputMemBlock_257 <= outputMemBlock_258;
    end
    if (nextBitValid) begin
      outputMemBlock_258 <= outputMemBlock_259;
    end
    if (nextBitValid) begin
      outputMemBlock_259 <= outputMemBlock_260;
    end
    if (nextBitValid) begin
      outputMemBlock_260 <= outputMemBlock_261;
    end
    if (nextBitValid) begin
      outputMemBlock_261 <= outputMemBlock_262;
    end
    if (nextBitValid) begin
      outputMemBlock_262 <= outputMemBlock_263;
    end
    if (nextBitValid) begin
      outputMemBlock_263 <= outputMemBlock_264;
    end
    if (nextBitValid) begin
      outputMemBlock_264 <= outputMemBlock_265;
    end
    if (nextBitValid) begin
      outputMemBlock_265 <= outputMemBlock_266;
    end
    if (nextBitValid) begin
      outputMemBlock_266 <= outputMemBlock_267;
    end
    if (nextBitValid) begin
      outputMemBlock_267 <= outputMemBlock_268;
    end
    if (nextBitValid) begin
      outputMemBlock_268 <= outputMemBlock_269;
    end
    if (nextBitValid) begin
      outputMemBlock_269 <= outputMemBlock_270;
    end
    if (nextBitValid) begin
      outputMemBlock_270 <= outputMemBlock_271;
    end
    if (nextBitValid) begin
      outputMemBlock_271 <= outputMemBlock_272;
    end
    if (nextBitValid) begin
      outputMemBlock_272 <= outputMemBlock_273;
    end
    if (nextBitValid) begin
      outputMemBlock_273 <= outputMemBlock_274;
    end
    if (nextBitValid) begin
      outputMemBlock_274 <= outputMemBlock_275;
    end
    if (nextBitValid) begin
      outputMemBlock_275 <= outputMemBlock_276;
    end
    if (nextBitValid) begin
      outputMemBlock_276 <= outputMemBlock_277;
    end
    if (nextBitValid) begin
      outputMemBlock_277 <= outputMemBlock_278;
    end
    if (nextBitValid) begin
      outputMemBlock_278 <= outputMemBlock_279;
    end
    if (nextBitValid) begin
      outputMemBlock_279 <= outputMemBlock_280;
    end
    if (nextBitValid) begin
      outputMemBlock_280 <= outputMemBlock_281;
    end
    if (nextBitValid) begin
      outputMemBlock_281 <= outputMemBlock_282;
    end
    if (nextBitValid) begin
      outputMemBlock_282 <= outputMemBlock_283;
    end
    if (nextBitValid) begin
      outputMemBlock_283 <= outputMemBlock_284;
    end
    if (nextBitValid) begin
      outputMemBlock_284 <= outputMemBlock_285;
    end
    if (nextBitValid) begin
      outputMemBlock_285 <= outputMemBlock_286;
    end
    if (nextBitValid) begin
      outputMemBlock_286 <= outputMemBlock_287;
    end
    if (nextBitValid) begin
      outputMemBlock_287 <= outputMemBlock_288;
    end
    if (nextBitValid) begin
      outputMemBlock_288 <= outputMemBlock_289;
    end
    if (nextBitValid) begin
      outputMemBlock_289 <= outputMemBlock_290;
    end
    if (nextBitValid) begin
      outputMemBlock_290 <= outputMemBlock_291;
    end
    if (nextBitValid) begin
      outputMemBlock_291 <= outputMemBlock_292;
    end
    if (nextBitValid) begin
      outputMemBlock_292 <= outputMemBlock_293;
    end
    if (nextBitValid) begin
      outputMemBlock_293 <= outputMemBlock_294;
    end
    if (nextBitValid) begin
      outputMemBlock_294 <= outputMemBlock_295;
    end
    if (nextBitValid) begin
      outputMemBlock_295 <= outputMemBlock_296;
    end
    if (nextBitValid) begin
      outputMemBlock_296 <= outputMemBlock_297;
    end
    if (nextBitValid) begin
      outputMemBlock_297 <= outputMemBlock_298;
    end
    if (nextBitValid) begin
      outputMemBlock_298 <= outputMemBlock_299;
    end
    if (nextBitValid) begin
      outputMemBlock_299 <= outputMemBlock_300;
    end
    if (nextBitValid) begin
      outputMemBlock_300 <= outputMemBlock_301;
    end
    if (nextBitValid) begin
      outputMemBlock_301 <= outputMemBlock_302;
    end
    if (nextBitValid) begin
      outputMemBlock_302 <= outputMemBlock_303;
    end
    if (nextBitValid) begin
      outputMemBlock_303 <= outputMemBlock_304;
    end
    if (nextBitValid) begin
      outputMemBlock_304 <= outputMemBlock_305;
    end
    if (nextBitValid) begin
      outputMemBlock_305 <= outputMemBlock_306;
    end
    if (nextBitValid) begin
      outputMemBlock_306 <= outputMemBlock_307;
    end
    if (nextBitValid) begin
      outputMemBlock_307 <= outputMemBlock_308;
    end
    if (nextBitValid) begin
      outputMemBlock_308 <= outputMemBlock_309;
    end
    if (nextBitValid) begin
      outputMemBlock_309 <= outputMemBlock_310;
    end
    if (nextBitValid) begin
      outputMemBlock_310 <= outputMemBlock_311;
    end
    if (nextBitValid) begin
      outputMemBlock_311 <= outputMemBlock_312;
    end
    if (nextBitValid) begin
      outputMemBlock_312 <= outputMemBlock_313;
    end
    if (nextBitValid) begin
      outputMemBlock_313 <= outputMemBlock_314;
    end
    if (nextBitValid) begin
      outputMemBlock_314 <= outputMemBlock_315;
    end
    if (nextBitValid) begin
      outputMemBlock_315 <= outputMemBlock_316;
    end
    if (nextBitValid) begin
      outputMemBlock_316 <= outputMemBlock_317;
    end
    if (nextBitValid) begin
      outputMemBlock_317 <= outputMemBlock_318;
    end
    if (nextBitValid) begin
      outputMemBlock_318 <= outputMemBlock_319;
    end
    if (nextBitValid) begin
      outputMemBlock_319 <= outputMemBlock_320;
    end
    if (nextBitValid) begin
      outputMemBlock_320 <= outputMemBlock_321;
    end
    if (nextBitValid) begin
      outputMemBlock_321 <= outputMemBlock_322;
    end
    if (nextBitValid) begin
      outputMemBlock_322 <= outputMemBlock_323;
    end
    if (nextBitValid) begin
      outputMemBlock_323 <= outputMemBlock_324;
    end
    if (nextBitValid) begin
      outputMemBlock_324 <= outputMemBlock_325;
    end
    if (nextBitValid) begin
      outputMemBlock_325 <= outputMemBlock_326;
    end
    if (nextBitValid) begin
      outputMemBlock_326 <= outputMemBlock_327;
    end
    if (nextBitValid) begin
      outputMemBlock_327 <= outputMemBlock_328;
    end
    if (nextBitValid) begin
      outputMemBlock_328 <= outputMemBlock_329;
    end
    if (nextBitValid) begin
      outputMemBlock_329 <= outputMemBlock_330;
    end
    if (nextBitValid) begin
      outputMemBlock_330 <= outputMemBlock_331;
    end
    if (nextBitValid) begin
      outputMemBlock_331 <= outputMemBlock_332;
    end
    if (nextBitValid) begin
      outputMemBlock_332 <= outputMemBlock_333;
    end
    if (nextBitValid) begin
      outputMemBlock_333 <= outputMemBlock_334;
    end
    if (nextBitValid) begin
      outputMemBlock_334 <= outputMemBlock_335;
    end
    if (nextBitValid) begin
      outputMemBlock_335 <= outputMemBlock_336;
    end
    if (nextBitValid) begin
      outputMemBlock_336 <= outputMemBlock_337;
    end
    if (nextBitValid) begin
      outputMemBlock_337 <= outputMemBlock_338;
    end
    if (nextBitValid) begin
      outputMemBlock_338 <= outputMemBlock_339;
    end
    if (nextBitValid) begin
      outputMemBlock_339 <= outputMemBlock_340;
    end
    if (nextBitValid) begin
      outputMemBlock_340 <= outputMemBlock_341;
    end
    if (nextBitValid) begin
      outputMemBlock_341 <= outputMemBlock_342;
    end
    if (nextBitValid) begin
      outputMemBlock_342 <= outputMemBlock_343;
    end
    if (nextBitValid) begin
      outputMemBlock_343 <= outputMemBlock_344;
    end
    if (nextBitValid) begin
      outputMemBlock_344 <= outputMemBlock_345;
    end
    if (nextBitValid) begin
      outputMemBlock_345 <= outputMemBlock_346;
    end
    if (nextBitValid) begin
      outputMemBlock_346 <= outputMemBlock_347;
    end
    if (nextBitValid) begin
      outputMemBlock_347 <= outputMemBlock_348;
    end
    if (nextBitValid) begin
      outputMemBlock_348 <= outputMemBlock_349;
    end
    if (nextBitValid) begin
      outputMemBlock_349 <= outputMemBlock_350;
    end
    if (nextBitValid) begin
      outputMemBlock_350 <= outputMemBlock_351;
    end
    if (nextBitValid) begin
      outputMemBlock_351 <= outputMemBlock_352;
    end
    if (nextBitValid) begin
      outputMemBlock_352 <= outputMemBlock_353;
    end
    if (nextBitValid) begin
      outputMemBlock_353 <= outputMemBlock_354;
    end
    if (nextBitValid) begin
      outputMemBlock_354 <= outputMemBlock_355;
    end
    if (nextBitValid) begin
      outputMemBlock_355 <= outputMemBlock_356;
    end
    if (nextBitValid) begin
      outputMemBlock_356 <= outputMemBlock_357;
    end
    if (nextBitValid) begin
      outputMemBlock_357 <= outputMemBlock_358;
    end
    if (nextBitValid) begin
      outputMemBlock_358 <= outputMemBlock_359;
    end
    if (nextBitValid) begin
      outputMemBlock_359 <= outputMemBlock_360;
    end
    if (nextBitValid) begin
      outputMemBlock_360 <= outputMemBlock_361;
    end
    if (nextBitValid) begin
      outputMemBlock_361 <= outputMemBlock_362;
    end
    if (nextBitValid) begin
      outputMemBlock_362 <= outputMemBlock_363;
    end
    if (nextBitValid) begin
      outputMemBlock_363 <= outputMemBlock_364;
    end
    if (nextBitValid) begin
      outputMemBlock_364 <= outputMemBlock_365;
    end
    if (nextBitValid) begin
      outputMemBlock_365 <= outputMemBlock_366;
    end
    if (nextBitValid) begin
      outputMemBlock_366 <= outputMemBlock_367;
    end
    if (nextBitValid) begin
      outputMemBlock_367 <= outputMemBlock_368;
    end
    if (nextBitValid) begin
      outputMemBlock_368 <= outputMemBlock_369;
    end
    if (nextBitValid) begin
      outputMemBlock_369 <= outputMemBlock_370;
    end
    if (nextBitValid) begin
      outputMemBlock_370 <= outputMemBlock_371;
    end
    if (nextBitValid) begin
      outputMemBlock_371 <= outputMemBlock_372;
    end
    if (nextBitValid) begin
      outputMemBlock_372 <= outputMemBlock_373;
    end
    if (nextBitValid) begin
      outputMemBlock_373 <= outputMemBlock_374;
    end
    if (nextBitValid) begin
      outputMemBlock_374 <= outputMemBlock_375;
    end
    if (nextBitValid) begin
      outputMemBlock_375 <= outputMemBlock_376;
    end
    if (nextBitValid) begin
      outputMemBlock_376 <= outputMemBlock_377;
    end
    if (nextBitValid) begin
      outputMemBlock_377 <= outputMemBlock_378;
    end
    if (nextBitValid) begin
      outputMemBlock_378 <= outputMemBlock_379;
    end
    if (nextBitValid) begin
      outputMemBlock_379 <= outputMemBlock_380;
    end
    if (nextBitValid) begin
      outputMemBlock_380 <= outputMemBlock_381;
    end
    if (nextBitValid) begin
      outputMemBlock_381 <= outputMemBlock_382;
    end
    if (nextBitValid) begin
      outputMemBlock_382 <= outputMemBlock_383;
    end
    if (nextBitValid) begin
      outputMemBlock_383 <= outputMemBlock_384;
    end
    if (nextBitValid) begin
      outputMemBlock_384 <= outputMemBlock_385;
    end
    if (nextBitValid) begin
      outputMemBlock_385 <= outputMemBlock_386;
    end
    if (nextBitValid) begin
      outputMemBlock_386 <= outputMemBlock_387;
    end
    if (nextBitValid) begin
      outputMemBlock_387 <= outputMemBlock_388;
    end
    if (nextBitValid) begin
      outputMemBlock_388 <= outputMemBlock_389;
    end
    if (nextBitValid) begin
      outputMemBlock_389 <= outputMemBlock_390;
    end
    if (nextBitValid) begin
      outputMemBlock_390 <= outputMemBlock_391;
    end
    if (nextBitValid) begin
      outputMemBlock_391 <= outputMemBlock_392;
    end
    if (nextBitValid) begin
      outputMemBlock_392 <= outputMemBlock_393;
    end
    if (nextBitValid) begin
      outputMemBlock_393 <= outputMemBlock_394;
    end
    if (nextBitValid) begin
      outputMemBlock_394 <= outputMemBlock_395;
    end
    if (nextBitValid) begin
      outputMemBlock_395 <= outputMemBlock_396;
    end
    if (nextBitValid) begin
      outputMemBlock_396 <= outputMemBlock_397;
    end
    if (nextBitValid) begin
      outputMemBlock_397 <= outputMemBlock_398;
    end
    if (nextBitValid) begin
      outputMemBlock_398 <= outputMemBlock_399;
    end
    if (nextBitValid) begin
      outputMemBlock_399 <= outputMemBlock_400;
    end
    if (nextBitValid) begin
      outputMemBlock_400 <= outputMemBlock_401;
    end
    if (nextBitValid) begin
      outputMemBlock_401 <= outputMemBlock_402;
    end
    if (nextBitValid) begin
      outputMemBlock_402 <= outputMemBlock_403;
    end
    if (nextBitValid) begin
      outputMemBlock_403 <= outputMemBlock_404;
    end
    if (nextBitValid) begin
      outputMemBlock_404 <= outputMemBlock_405;
    end
    if (nextBitValid) begin
      outputMemBlock_405 <= outputMemBlock_406;
    end
    if (nextBitValid) begin
      outputMemBlock_406 <= outputMemBlock_407;
    end
    if (nextBitValid) begin
      outputMemBlock_407 <= outputMemBlock_408;
    end
    if (nextBitValid) begin
      outputMemBlock_408 <= outputMemBlock_409;
    end
    if (nextBitValid) begin
      outputMemBlock_409 <= outputMemBlock_410;
    end
    if (nextBitValid) begin
      outputMemBlock_410 <= outputMemBlock_411;
    end
    if (nextBitValid) begin
      outputMemBlock_411 <= outputMemBlock_412;
    end
    if (nextBitValid) begin
      outputMemBlock_412 <= outputMemBlock_413;
    end
    if (nextBitValid) begin
      outputMemBlock_413 <= outputMemBlock_414;
    end
    if (nextBitValid) begin
      outputMemBlock_414 <= outputMemBlock_415;
    end
    if (nextBitValid) begin
      outputMemBlock_415 <= outputMemBlock_416;
    end
    if (nextBitValid) begin
      outputMemBlock_416 <= outputMemBlock_417;
    end
    if (nextBitValid) begin
      outputMemBlock_417 <= outputMemBlock_418;
    end
    if (nextBitValid) begin
      outputMemBlock_418 <= outputMemBlock_419;
    end
    if (nextBitValid) begin
      outputMemBlock_419 <= outputMemBlock_420;
    end
    if (nextBitValid) begin
      outputMemBlock_420 <= outputMemBlock_421;
    end
    if (nextBitValid) begin
      outputMemBlock_421 <= outputMemBlock_422;
    end
    if (nextBitValid) begin
      outputMemBlock_422 <= outputMemBlock_423;
    end
    if (nextBitValid) begin
      outputMemBlock_423 <= outputMemBlock_424;
    end
    if (nextBitValid) begin
      outputMemBlock_424 <= outputMemBlock_425;
    end
    if (nextBitValid) begin
      outputMemBlock_425 <= outputMemBlock_426;
    end
    if (nextBitValid) begin
      outputMemBlock_426 <= outputMemBlock_427;
    end
    if (nextBitValid) begin
      outputMemBlock_427 <= outputMemBlock_428;
    end
    if (nextBitValid) begin
      outputMemBlock_428 <= outputMemBlock_429;
    end
    if (nextBitValid) begin
      outputMemBlock_429 <= outputMemBlock_430;
    end
    if (nextBitValid) begin
      outputMemBlock_430 <= outputMemBlock_431;
    end
    if (nextBitValid) begin
      outputMemBlock_431 <= outputMemBlock_432;
    end
    if (nextBitValid) begin
      outputMemBlock_432 <= outputMemBlock_433;
    end
    if (nextBitValid) begin
      outputMemBlock_433 <= outputMemBlock_434;
    end
    if (nextBitValid) begin
      outputMemBlock_434 <= outputMemBlock_435;
    end
    if (nextBitValid) begin
      outputMemBlock_435 <= outputMemBlock_436;
    end
    if (nextBitValid) begin
      outputMemBlock_436 <= outputMemBlock_437;
    end
    if (nextBitValid) begin
      outputMemBlock_437 <= outputMemBlock_438;
    end
    if (nextBitValid) begin
      outputMemBlock_438 <= outputMemBlock_439;
    end
    if (nextBitValid) begin
      outputMemBlock_439 <= outputMemBlock_440;
    end
    if (nextBitValid) begin
      outputMemBlock_440 <= outputMemBlock_441;
    end
    if (nextBitValid) begin
      outputMemBlock_441 <= outputMemBlock_442;
    end
    if (nextBitValid) begin
      outputMemBlock_442 <= outputMemBlock_443;
    end
    if (nextBitValid) begin
      outputMemBlock_443 <= outputMemBlock_444;
    end
    if (nextBitValid) begin
      outputMemBlock_444 <= outputMemBlock_445;
    end
    if (nextBitValid) begin
      outputMemBlock_445 <= outputMemBlock_446;
    end
    if (nextBitValid) begin
      outputMemBlock_446 <= outputMemBlock_447;
    end
    if (nextBitValid) begin
      outputMemBlock_447 <= outputMemBlock_448;
    end
    if (nextBitValid) begin
      outputMemBlock_448 <= outputMemBlock_449;
    end
    if (nextBitValid) begin
      outputMemBlock_449 <= outputMemBlock_450;
    end
    if (nextBitValid) begin
      outputMemBlock_450 <= outputMemBlock_451;
    end
    if (nextBitValid) begin
      outputMemBlock_451 <= outputMemBlock_452;
    end
    if (nextBitValid) begin
      outputMemBlock_452 <= outputMemBlock_453;
    end
    if (nextBitValid) begin
      outputMemBlock_453 <= outputMemBlock_454;
    end
    if (nextBitValid) begin
      outputMemBlock_454 <= outputMemBlock_455;
    end
    if (nextBitValid) begin
      outputMemBlock_455 <= outputMemBlock_456;
    end
    if (nextBitValid) begin
      outputMemBlock_456 <= outputMemBlock_457;
    end
    if (nextBitValid) begin
      outputMemBlock_457 <= outputMemBlock_458;
    end
    if (nextBitValid) begin
      outputMemBlock_458 <= outputMemBlock_459;
    end
    if (nextBitValid) begin
      outputMemBlock_459 <= outputMemBlock_460;
    end
    if (nextBitValid) begin
      outputMemBlock_460 <= outputMemBlock_461;
    end
    if (nextBitValid) begin
      outputMemBlock_461 <= outputMemBlock_462;
    end
    if (nextBitValid) begin
      outputMemBlock_462 <= outputMemBlock_463;
    end
    if (nextBitValid) begin
      outputMemBlock_463 <= outputMemBlock_464;
    end
    if (nextBitValid) begin
      outputMemBlock_464 <= outputMemBlock_465;
    end
    if (nextBitValid) begin
      outputMemBlock_465 <= outputMemBlock_466;
    end
    if (nextBitValid) begin
      outputMemBlock_466 <= outputMemBlock_467;
    end
    if (nextBitValid) begin
      outputMemBlock_467 <= outputMemBlock_468;
    end
    if (nextBitValid) begin
      outputMemBlock_468 <= outputMemBlock_469;
    end
    if (nextBitValid) begin
      outputMemBlock_469 <= outputMemBlock_470;
    end
    if (nextBitValid) begin
      outputMemBlock_470 <= outputMemBlock_471;
    end
    if (nextBitValid) begin
      outputMemBlock_471 <= outputMemBlock_472;
    end
    if (nextBitValid) begin
      outputMemBlock_472 <= outputMemBlock_473;
    end
    if (nextBitValid) begin
      outputMemBlock_473 <= outputMemBlock_474;
    end
    if (nextBitValid) begin
      outputMemBlock_474 <= outputMemBlock_475;
    end
    if (nextBitValid) begin
      outputMemBlock_475 <= outputMemBlock_476;
    end
    if (nextBitValid) begin
      outputMemBlock_476 <= outputMemBlock_477;
    end
    if (nextBitValid) begin
      outputMemBlock_477 <= outputMemBlock_478;
    end
    if (nextBitValid) begin
      outputMemBlock_478 <= outputMemBlock_479;
    end
    if (nextBitValid) begin
      outputMemBlock_479 <= outputMemBlock_480;
    end
    if (nextBitValid) begin
      outputMemBlock_480 <= outputMemBlock_481;
    end
    if (nextBitValid) begin
      outputMemBlock_481 <= outputMemBlock_482;
    end
    if (nextBitValid) begin
      outputMemBlock_482 <= outputMemBlock_483;
    end
    if (nextBitValid) begin
      outputMemBlock_483 <= outputMemBlock_484;
    end
    if (nextBitValid) begin
      outputMemBlock_484 <= outputMemBlock_485;
    end
    if (nextBitValid) begin
      outputMemBlock_485 <= outputMemBlock_486;
    end
    if (nextBitValid) begin
      outputMemBlock_486 <= outputMemBlock_487;
    end
    if (nextBitValid) begin
      outputMemBlock_487 <= outputMemBlock_488;
    end
    if (nextBitValid) begin
      outputMemBlock_488 <= outputMemBlock_489;
    end
    if (nextBitValid) begin
      outputMemBlock_489 <= outputMemBlock_490;
    end
    if (nextBitValid) begin
      outputMemBlock_490 <= outputMemBlock_491;
    end
    if (nextBitValid) begin
      outputMemBlock_491 <= outputMemBlock_492;
    end
    if (nextBitValid) begin
      outputMemBlock_492 <= outputMemBlock_493;
    end
    if (nextBitValid) begin
      outputMemBlock_493 <= outputMemBlock_494;
    end
    if (nextBitValid) begin
      outputMemBlock_494 <= outputMemBlock_495;
    end
    if (nextBitValid) begin
      outputMemBlock_495 <= outputMemBlock_496;
    end
    if (nextBitValid) begin
      outputMemBlock_496 <= outputMemBlock_497;
    end
    if (nextBitValid) begin
      outputMemBlock_497 <= outputMemBlock_498;
    end
    if (nextBitValid) begin
      outputMemBlock_498 <= outputMemBlock_499;
    end
    if (nextBitValid) begin
      outputMemBlock_499 <= outputMemBlock_500;
    end
    if (nextBitValid) begin
      outputMemBlock_500 <= outputMemBlock_501;
    end
    if (nextBitValid) begin
      outputMemBlock_501 <= outputMemBlock_502;
    end
    if (nextBitValid) begin
      outputMemBlock_502 <= outputMemBlock_503;
    end
    if (nextBitValid) begin
      outputMemBlock_503 <= outputMemBlock_504;
    end
    if (nextBitValid) begin
      outputMemBlock_504 <= outputMemBlock_505;
    end
    if (nextBitValid) begin
      outputMemBlock_505 <= outputMemBlock_506;
    end
    if (nextBitValid) begin
      outputMemBlock_506 <= outputMemBlock_507;
    end
    if (nextBitValid) begin
      outputMemBlock_507 <= outputMemBlock_508;
    end
    if (nextBitValid) begin
      outputMemBlock_508 <= outputMemBlock_509;
    end
    if (nextBitValid) begin
      outputMemBlock_509 <= outputMemBlock_510;
    end
    if (nextBitValid) begin
      outputMemBlock_510 <= outputMemBlock_511;
    end
    if (nextBitValid) begin
      outputMemBlock_511 <= nextBit;
    end
    if (reset) begin
      outputBits <= 10'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputBits <= 10'h0;
      end else begin
        if (nextBitValid) begin
          outputBits <= _T_1588;
        end
      end
    end
  end
endmodule
module StreamingCore(
  input   clock,
  input   reset,
  output [63:0] io_inputMemAddr,
  output  io_inputMemAddrValid,
  input   io_inputMemAddrReady,
  input  [511:0] io_inputMemBlock,
  input   io_inputMemBlockValid,
  output  io_inputMemBlockReady,
  output [63:0] io_outputMemAddr,
  output  io_outputMemAddrValid,
  input   io_outputMemAddrReady,
  output [511:0] io_outputMemBlock,
  output  io_outputMemBlockValid,
  input   io_outputMemBlockReady,
  output  io_inputFinished,
  output  io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [511:0] core_io_inputMemBlock;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [511:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _GEN_26;
  reg  initDone;
  reg [31:0] _GEN_27;
  reg [63:0] inputBitsRemaining;
  reg [63:0] _GEN_28;
  reg  coreInputFinished;
  reg [31:0] _GEN_29;
  reg [63:0] outputBits;
  reg [63:0] _GEN_30;
  reg  outputLengthCommitted;
  reg [31:0] _GEN_31;
  reg [63:0] inputMemAddr;
  reg [63:0] _GEN_32;
  reg [63:0] outputMemAddr;
  reg [63:0] _GEN_33;
  reg [63:0] outputLenAddr;
  reg [63:0] _GEN_34;
  reg  outputMemFlushed;
  reg [31:0] _GEN_35;
  reg  inputAddressAccepted;
  reg [31:0] _GEN_36;
  wire  _T_42;
  wire  _T_43;
  wire  _T_45;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_51;
  wire  _GEN_0;
  wire  inputBlockReadable;
  wire  _T_54;
  wire  _T_55;
  wire  _T_57;
  wire [9:0] _T_59;
  wire [9:0] _T_60;
  wire [63:0] _T_61;
  wire [63:0] _T_62;
  wire [63:0] _T_63;
  wire [64:0] _T_65;
  wire [63:0] _T_66;
  wire [63:0] _GEN_1;
  wire [63:0] _GEN_2;
  wire [63:0] _GEN_3;
  wire [63:0] _GEN_4;
  wire  _GEN_5;
  wire  _GEN_6;
  wire  _T_71;
  wire [64:0] _T_75;
  wire [63:0] _T_76;
  wire [63:0] _T_78;
  wire [64:0] _T_80;
  wire [63:0] _T_81;
  wire [63:0] _GEN_7;
  wire [63:0] _GEN_8;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _T_87;
  wire  _GEN_16;
  reg  outputAddressAccepted;
  reg [31:0] _GEN_37;
  wire [63:0] _T_90;
  wire  _T_92;
  wire  _T_94;
  wire  _T_95;
  wire  _T_96;
  wire  _T_97;
  wire  _T_98;
  wire  _GEN_17;
  wire [511:0] _T_100;
  wire  _T_101;
  wire  _GEN_18;
  wire  _T_106;
  wire [63:0] _GEN_25;
  wire [64:0] _T_107;
  wire [63:0] _T_108;
  wire [64:0] _T_110;
  wire [63:0] _T_111;
  wire [63:0] _GEN_19;
  wire [63:0] _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemAddrValid = _T_50;
  assign io_inputMemBlockReady = inputAddressAccepted;
  assign io_outputMemAddr = _T_90;
  assign io_outputMemAddrValid = _T_97;
  assign io_outputMemBlock = _T_100;
  assign io_outputMemBlockValid = outputAddressAccepted;
  assign io_inputFinished = _T_45;
  assign io_outputFinished = outputLengthCommitted;
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemBlockValid = _T_55;
  assign core_io_inputBits = _T_60;
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemFlushed = _T_101;
  assign _T_42 = inputAddressAccepted == 1'h0;
  assign _T_43 = initDone & core_io_inputMemConsumed;
  assign _T_45 = inputBitsRemaining == 64'h0;
  assign _T_47 = _T_45 == 1'h0;
  assign _T_48 = _T_43 & _T_47;
  assign _T_49 = isInit | _T_48;
  assign _T_50 = _T_42 & _T_49;
  assign _T_51 = io_inputMemAddrValid & io_inputMemAddrReady;
  assign _GEN_0 = _T_51 ? 1'h1 : inputAddressAccepted;
  assign inputBlockReadable = _T_54;
  assign _T_54 = inputAddressAccepted & io_inputMemBlockValid;
  assign _T_55 = inputBlockReadable & initDone;
  assign _T_57 = inputBitsRemaining > 64'h200;
  assign _T_59 = inputBitsRemaining[9:0];
  assign _T_60 = _T_57 ? 10'h200 : _T_59;
  assign _T_61 = io_inputMemBlock[63:0];
  assign _T_62 = io_inputMemBlock[127:64];
  assign _T_63 = io_inputMemBlock[191:128];
  assign _T_65 = _T_63 + 64'h40;
  assign _T_66 = _T_65[63:0];
  assign _GEN_1 = isInit ? _T_61 : inputMemAddr;
  assign _GEN_2 = isInit ? _T_62 : inputBitsRemaining;
  assign _GEN_3 = isInit ? _T_66 : outputMemAddr;
  assign _GEN_4 = isInit ? _T_63 : outputLenAddr;
  assign _GEN_5 = isInit ? 1'h0 : isInit;
  assign _GEN_6 = isInit ? 1'h1 : initDone;
  assign _T_71 = isInit == 1'h0;
  assign _T_75 = inputBitsRemaining - 64'h200;
  assign _T_76 = _T_75[63:0];
  assign _T_78 = _T_57 ? _T_76 : 64'h0;
  assign _T_80 = inputMemAddr + 64'h40;
  assign _T_81 = _T_80[63:0];
  assign _GEN_7 = _T_71 ? _T_78 : _GEN_2;
  assign _GEN_8 = _T_71 ? _T_81 : _GEN_1;
  assign _GEN_9 = inputBlockReadable ? _GEN_8 : inputMemAddr;
  assign _GEN_10 = inputBlockReadable ? _GEN_7 : inputBitsRemaining;
  assign _GEN_11 = inputBlockReadable ? _GEN_3 : outputMemAddr;
  assign _GEN_12 = inputBlockReadable ? _GEN_4 : outputLenAddr;
  assign _GEN_13 = inputBlockReadable ? _GEN_5 : isInit;
  assign _GEN_14 = inputBlockReadable ? _GEN_6 : initDone;
  assign _GEN_15 = inputBlockReadable ? 1'h0 : _GEN_0;
  assign _T_87 = core_io_inputMemConsumed & _T_45;
  assign _GEN_16 = _T_87 ? 1'h1 : coreInputFinished;
  assign _T_90 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_92 = outputAddressAccepted == 1'h0;
  assign _T_94 = outputLengthCommitted == 1'h0;
  assign _T_95 = core_io_outputFinished & _T_94;
  assign _T_96 = core_io_outputMemBlockValid | _T_95;
  assign _T_97 = _T_92 & _T_96;
  assign _T_98 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_17 = _T_98 ? 1'h1 : outputAddressAccepted;
  assign _T_100 = core_io_outputFinished ? {{448'd0}, outputBits} : core_io_outputMemBlock;
  assign _T_101 = outputAddressAccepted & io_outputMemBlockReady;
  assign _GEN_18 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _T_106 = core_io_outputFinished == 1'h0;
  assign _GEN_25 = {{54'd0}, core_io_outputBits};
  assign _T_107 = outputBits + _GEN_25;
  assign _T_108 = _T_107[63:0];
  assign _T_110 = outputMemAddr + 64'h40;
  assign _T_111 = _T_110[63:0];
  assign _GEN_19 = _T_106 ? _T_108 : outputBits;
  assign _GEN_20 = _T_106 ? _T_111 : _GEN_11;
  assign _GEN_21 = _T_101 ? 1'h0 : _GEN_17;
  assign _GEN_22 = _T_101 ? _GEN_18 : outputLengthCommitted;
  assign _GEN_23 = _T_101 ? _GEN_19 : outputBits;
  assign _GEN_24 = _T_101 ? _GEN_20 : _GEN_11;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_26 = {1{$random}};
  isInit = _GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_27 = {1{$random}};
  initDone = _GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_28 = {2{$random}};
  inputBitsRemaining = _GEN_28[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_29 = {1{$random}};
  coreInputFinished = _GEN_29[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_30 = {2{$random}};
  outputBits = _GEN_30[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_31 = {1{$random}};
  outputLengthCommitted = _GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_32 = {2{$random}};
  inputMemAddr = _GEN_32[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_33 = {2{$random}};
  outputMemAddr = _GEN_33[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_34 = {2{$random}};
  outputLenAddr = _GEN_34[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_35 = {1{$random}};
  outputMemFlushed = _GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_36 = {1{$random}};
  inputAddressAccepted = _GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_37 = {1{$random}};
  outputAddressAccepted = _GEN_37[0:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          isInit <= 1'h0;
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          initDone <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 64'h1;
    end else begin
      if (inputBlockReadable) begin
        if (_T_71) begin
          if (_T_57) begin
            inputBitsRemaining <= _T_76;
          end else begin
            inputBitsRemaining <= 64'h0;
          end
        end else begin
          if (isInit) begin
            inputBitsRemaining <= _T_62;
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_87) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 64'h0;
    end else begin
      if (_T_101) begin
        if (_T_106) begin
          outputBits <= _T_108;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_101) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 64'h0;
    end else begin
      if (inputBlockReadable) begin
        if (_T_71) begin
          inputMemAddr <= _T_81;
        end else begin
          if (isInit) begin
            inputMemAddr <= _T_61;
          end
        end
      end
    end
    if (_T_101) begin
      if (_T_106) begin
        outputMemAddr <= _T_111;
      end else begin
        if (inputBlockReadable) begin
          if (isInit) begin
            outputMemAddr <= _T_66;
          end
        end
      end
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          outputMemAddr <= _T_66;
        end
      end
    end
    if (inputBlockReadable) begin
      if (isInit) begin
        outputLenAddr <= _T_63;
      end
    end
    if (reset) begin
      outputMemFlushed <= 1'h0;
    end
    if (reset) begin
      inputAddressAccepted <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        inputAddressAccepted <= 1'h0;
      end else begin
        if (_T_51) begin
          inputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_101) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_98) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
  end
endmodule
module StreamingCore_1(
  input   clock,
  input   reset,
  output [63:0] io_inputMemAddr,
  output  io_inputMemAddrValid,
  input   io_inputMemAddrReady,
  input  [511:0] io_inputMemBlock,
  input   io_inputMemBlockValid,
  output  io_inputMemBlockReady,
  output [63:0] io_outputMemAddr,
  output  io_outputMemAddrValid,
  input   io_outputMemAddrReady,
  output [511:0] io_outputMemBlock,
  output  io_outputMemBlockValid,
  input   io_outputMemBlockReady,
  output  io_inputFinished,
  output  io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [511:0] core_io_inputMemBlock;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [511:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _GEN_26;
  reg  initDone;
  reg [31:0] _GEN_27;
  reg [63:0] inputBitsRemaining;
  reg [63:0] _GEN_28;
  reg  coreInputFinished;
  reg [31:0] _GEN_29;
  reg [63:0] outputBits;
  reg [63:0] _GEN_30;
  reg  outputLengthCommitted;
  reg [31:0] _GEN_31;
  reg [63:0] inputMemAddr;
  reg [63:0] _GEN_32;
  reg [63:0] outputMemAddr;
  reg [63:0] _GEN_33;
  reg [63:0] outputLenAddr;
  reg [63:0] _GEN_34;
  reg  outputMemFlushed;
  reg [31:0] _GEN_35;
  reg  inputAddressAccepted;
  reg [31:0] _GEN_36;
  wire  _T_42;
  wire  _T_43;
  wire  _T_45;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_51;
  wire  _GEN_0;
  wire  inputBlockReadable;
  wire  _T_54;
  wire  _T_55;
  wire  _T_57;
  wire [9:0] _T_59;
  wire [9:0] _T_60;
  wire [63:0] _T_61;
  wire [63:0] _T_62;
  wire [63:0] _T_63;
  wire [64:0] _T_65;
  wire [63:0] _T_66;
  wire [63:0] _GEN_1;
  wire [63:0] _GEN_2;
  wire [63:0] _GEN_3;
  wire [63:0] _GEN_4;
  wire  _GEN_5;
  wire  _GEN_6;
  wire  _T_71;
  wire [64:0] _T_75;
  wire [63:0] _T_76;
  wire [63:0] _T_78;
  wire [64:0] _T_80;
  wire [63:0] _T_81;
  wire [63:0] _GEN_7;
  wire [63:0] _GEN_8;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _T_87;
  wire  _GEN_16;
  reg  outputAddressAccepted;
  reg [31:0] _GEN_37;
  wire [63:0] _T_90;
  wire  _T_92;
  wire  _T_94;
  wire  _T_95;
  wire  _T_96;
  wire  _T_97;
  wire  _T_98;
  wire  _GEN_17;
  wire [511:0] _T_100;
  wire  _T_101;
  wire  _GEN_18;
  wire  _T_106;
  wire [63:0] _GEN_25;
  wire [64:0] _T_107;
  wire [63:0] _T_108;
  wire [64:0] _T_110;
  wire [63:0] _T_111;
  wire [63:0] _GEN_19;
  wire [63:0] _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemAddrValid = _T_50;
  assign io_inputMemBlockReady = inputAddressAccepted;
  assign io_outputMemAddr = _T_90;
  assign io_outputMemAddrValid = _T_97;
  assign io_outputMemBlock = _T_100;
  assign io_outputMemBlockValid = outputAddressAccepted;
  assign io_inputFinished = _T_45;
  assign io_outputFinished = outputLengthCommitted;
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemBlockValid = _T_55;
  assign core_io_inputBits = _T_60;
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemFlushed = _T_101;
  assign _T_42 = inputAddressAccepted == 1'h0;
  assign _T_43 = initDone & core_io_inputMemConsumed;
  assign _T_45 = inputBitsRemaining == 64'h0;
  assign _T_47 = _T_45 == 1'h0;
  assign _T_48 = _T_43 & _T_47;
  assign _T_49 = isInit | _T_48;
  assign _T_50 = _T_42 & _T_49;
  assign _T_51 = io_inputMemAddrValid & io_inputMemAddrReady;
  assign _GEN_0 = _T_51 ? 1'h1 : inputAddressAccepted;
  assign inputBlockReadable = _T_54;
  assign _T_54 = inputAddressAccepted & io_inputMemBlockValid;
  assign _T_55 = inputBlockReadable & initDone;
  assign _T_57 = inputBitsRemaining > 64'h200;
  assign _T_59 = inputBitsRemaining[9:0];
  assign _T_60 = _T_57 ? 10'h200 : _T_59;
  assign _T_61 = io_inputMemBlock[63:0];
  assign _T_62 = io_inputMemBlock[127:64];
  assign _T_63 = io_inputMemBlock[191:128];
  assign _T_65 = _T_63 + 64'h40;
  assign _T_66 = _T_65[63:0];
  assign _GEN_1 = isInit ? _T_61 : inputMemAddr;
  assign _GEN_2 = isInit ? _T_62 : inputBitsRemaining;
  assign _GEN_3 = isInit ? _T_66 : outputMemAddr;
  assign _GEN_4 = isInit ? _T_63 : outputLenAddr;
  assign _GEN_5 = isInit ? 1'h0 : isInit;
  assign _GEN_6 = isInit ? 1'h1 : initDone;
  assign _T_71 = isInit == 1'h0;
  assign _T_75 = inputBitsRemaining - 64'h200;
  assign _T_76 = _T_75[63:0];
  assign _T_78 = _T_57 ? _T_76 : 64'h0;
  assign _T_80 = inputMemAddr + 64'h40;
  assign _T_81 = _T_80[63:0];
  assign _GEN_7 = _T_71 ? _T_78 : _GEN_2;
  assign _GEN_8 = _T_71 ? _T_81 : _GEN_1;
  assign _GEN_9 = inputBlockReadable ? _GEN_8 : inputMemAddr;
  assign _GEN_10 = inputBlockReadable ? _GEN_7 : inputBitsRemaining;
  assign _GEN_11 = inputBlockReadable ? _GEN_3 : outputMemAddr;
  assign _GEN_12 = inputBlockReadable ? _GEN_4 : outputLenAddr;
  assign _GEN_13 = inputBlockReadable ? _GEN_5 : isInit;
  assign _GEN_14 = inputBlockReadable ? _GEN_6 : initDone;
  assign _GEN_15 = inputBlockReadable ? 1'h0 : _GEN_0;
  assign _T_87 = core_io_inputMemConsumed & _T_45;
  assign _GEN_16 = _T_87 ? 1'h1 : coreInputFinished;
  assign _T_90 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_92 = outputAddressAccepted == 1'h0;
  assign _T_94 = outputLengthCommitted == 1'h0;
  assign _T_95 = core_io_outputFinished & _T_94;
  assign _T_96 = core_io_outputMemBlockValid | _T_95;
  assign _T_97 = _T_92 & _T_96;
  assign _T_98 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_17 = _T_98 ? 1'h1 : outputAddressAccepted;
  assign _T_100 = core_io_outputFinished ? {{448'd0}, outputBits} : core_io_outputMemBlock;
  assign _T_101 = outputAddressAccepted & io_outputMemBlockReady;
  assign _GEN_18 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _T_106 = core_io_outputFinished == 1'h0;
  assign _GEN_25 = {{54'd0}, core_io_outputBits};
  assign _T_107 = outputBits + _GEN_25;
  assign _T_108 = _T_107[63:0];
  assign _T_110 = outputMemAddr + 64'h40;
  assign _T_111 = _T_110[63:0];
  assign _GEN_19 = _T_106 ? _T_108 : outputBits;
  assign _GEN_20 = _T_106 ? _T_111 : _GEN_11;
  assign _GEN_21 = _T_101 ? 1'h0 : _GEN_17;
  assign _GEN_22 = _T_101 ? _GEN_18 : outputLengthCommitted;
  assign _GEN_23 = _T_101 ? _GEN_19 : outputBits;
  assign _GEN_24 = _T_101 ? _GEN_20 : _GEN_11;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_26 = {1{$random}};
  isInit = _GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_27 = {1{$random}};
  initDone = _GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_28 = {2{$random}};
  inputBitsRemaining = _GEN_28[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_29 = {1{$random}};
  coreInputFinished = _GEN_29[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_30 = {2{$random}};
  outputBits = _GEN_30[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_31 = {1{$random}};
  outputLengthCommitted = _GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_32 = {2{$random}};
  inputMemAddr = _GEN_32[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_33 = {2{$random}};
  outputMemAddr = _GEN_33[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_34 = {2{$random}};
  outputLenAddr = _GEN_34[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_35 = {1{$random}};
  outputMemFlushed = _GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_36 = {1{$random}};
  inputAddressAccepted = _GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_37 = {1{$random}};
  outputAddressAccepted = _GEN_37[0:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          isInit <= 1'h0;
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          initDone <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 64'h1;
    end else begin
      if (inputBlockReadable) begin
        if (_T_71) begin
          if (_T_57) begin
            inputBitsRemaining <= _T_76;
          end else begin
            inputBitsRemaining <= 64'h0;
          end
        end else begin
          if (isInit) begin
            inputBitsRemaining <= _T_62;
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_87) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 64'h0;
    end else begin
      if (_T_101) begin
        if (_T_106) begin
          outputBits <= _T_108;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_101) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 64'h400000000;
    end else begin
      if (inputBlockReadable) begin
        if (_T_71) begin
          inputMemAddr <= _T_81;
        end else begin
          if (isInit) begin
            inputMemAddr <= _T_61;
          end
        end
      end
    end
    if (_T_101) begin
      if (_T_106) begin
        outputMemAddr <= _T_111;
      end else begin
        if (inputBlockReadable) begin
          if (isInit) begin
            outputMemAddr <= _T_66;
          end
        end
      end
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          outputMemAddr <= _T_66;
        end
      end
    end
    if (inputBlockReadable) begin
      if (isInit) begin
        outputLenAddr <= _T_63;
      end
    end
    if (reset) begin
      outputMemFlushed <= 1'h0;
    end
    if (reset) begin
      inputAddressAccepted <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        inputAddressAccepted <= 1'h0;
      end else begin
        if (_T_51) begin
          inputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_101) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_98) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
  end
endmodule
module StreamingWrapper(
  input   clock,
  input   reset,
  output [63:0] io_inputMemAddrs_0,
  output [63:0] io_inputMemAddrs_1,
  output  io_inputMemAddrValids_0,
  output  io_inputMemAddrValids_1,
  input   io_inputMemAddrReadys_0,
  input   io_inputMemAddrReadys_1,
  input  [511:0] io_inputMemBlocks_0,
  input  [511:0] io_inputMemBlocks_1,
  input   io_inputMemBlockValids_0,
  input   io_inputMemBlockValids_1,
  output  io_inputMemBlockReadys_0,
  output  io_inputMemBlockReadys_1,
  output [63:0] io_outputMemAddrs_0,
  output [63:0] io_outputMemAddrs_1,
  output  io_outputMemAddrValids_0,
  output  io_outputMemAddrValids_1,
  input   io_outputMemAddrReadys_0,
  input   io_outputMemAddrReadys_1,
  output [511:0] io_outputMemBlocks_0,
  output [511:0] io_outputMemBlocks_1,
  output  io_outputMemBlockValids_0,
  output  io_outputMemBlockValids_1,
  input   io_outputMemBlockReadys_0,
  input   io_outputMemBlockReadys_1,
  output  io_finished
);
  wire  StreamingCore_clock;
  wire  StreamingCore_reset;
  wire [63:0] StreamingCore_io_inputMemAddr;
  wire  StreamingCore_io_inputMemAddrValid;
  wire  StreamingCore_io_inputMemAddrReady;
  wire [511:0] StreamingCore_io_inputMemBlock;
  wire  StreamingCore_io_inputMemBlockValid;
  wire  StreamingCore_io_inputMemBlockReady;
  wire [63:0] StreamingCore_io_outputMemAddr;
  wire  StreamingCore_io_outputMemAddrValid;
  wire  StreamingCore_io_outputMemAddrReady;
  wire [511:0] StreamingCore_io_outputMemBlock;
  wire  StreamingCore_io_outputMemBlockValid;
  wire  StreamingCore_io_outputMemBlockReady;
  wire  StreamingCore_io_inputFinished;
  wire  StreamingCore_io_outputFinished;
  wire  StreamingCore_1_clock;
  wire  StreamingCore_1_reset;
  wire [63:0] StreamingCore_1_io_inputMemAddr;
  wire  StreamingCore_1_io_inputMemAddrValid;
  wire  StreamingCore_1_io_inputMemAddrReady;
  wire [511:0] StreamingCore_1_io_inputMemBlock;
  wire  StreamingCore_1_io_inputMemBlockValid;
  wire  StreamingCore_1_io_inputMemBlockReady;
  wire [63:0] StreamingCore_1_io_outputMemAddr;
  wire  StreamingCore_1_io_outputMemAddrValid;
  wire  StreamingCore_1_io_outputMemAddrReady;
  wire [511:0] StreamingCore_1_io_outputMemBlock;
  wire  StreamingCore_1_io_outputMemBlockValid;
  wire  StreamingCore_1_io_outputMemBlockReady;
  wire  StreamingCore_1_io_inputFinished;
  wire  StreamingCore_1_io_outputFinished;
  wire [63:0] cores_0_inputMemAddr;
  wire  cores_0_inputMemAddrValid;
  wire  cores_0_inputMemAddrReady;
  wire [511:0] cores_0_inputMemBlock;
  wire  cores_0_inputMemBlockValid;
  wire  cores_0_inputMemBlockReady;
  wire [63:0] cores_0_outputMemAddr;
  wire  cores_0_outputMemAddrValid;
  wire  cores_0_outputMemAddrReady;
  wire [511:0] cores_0_outputMemBlock;
  wire  cores_0_outputMemBlockValid;
  wire  cores_0_outputMemBlockReady;
  wire  cores_0_inputFinished;
  wire  cores_0_outputFinished;
  wire [63:0] cores_1_inputMemAddr;
  wire  cores_1_inputMemAddrValid;
  wire  cores_1_inputMemAddrReady;
  wire [511:0] cores_1_inputMemBlock;
  wire  cores_1_inputMemBlockValid;
  wire  cores_1_inputMemBlockReady;
  wire [63:0] cores_1_outputMemAddr;
  wire  cores_1_outputMemAddrValid;
  wire  cores_1_outputMemAddrReady;
  wire [511:0] cores_1_outputMemBlock;
  wire  cores_1_outputMemBlockValid;
  wire  cores_1_outputMemBlockReady;
  wire  cores_1_inputFinished;
  wire  cores_1_outputFinished;
  reg  _T_533;
  reg [31:0] _GEN_0;
  reg  _T_535;
  reg [31:0] _GEN_1;
  reg  _T_537;
  reg [31:0] _GEN_2;
  reg  _T_539;
  reg [31:0] _GEN_3;
  wire [63:0] _GEN_0_inputMemAddr;
  wire  _GEN_0_inputMemAddrValid;
  wire  _GEN_0_inputMemAddrReady;
  wire [511:0] _GEN_0_inputMemBlock;
  wire  _GEN_0_inputMemBlockValid;
  wire  _GEN_0_inputMemBlockReady;
  wire [63:0] _GEN_0_outputMemAddr;
  wire  _GEN_0_outputMemAddrValid;
  wire  _GEN_0_outputMemAddrReady;
  wire [511:0] _GEN_0_outputMemBlock;
  wire  _GEN_0_outputMemBlockValid;
  wire  _GEN_0_outputMemBlockReady;
  wire  _GEN_0_inputFinished;
  wire  _GEN_0_outputFinished;
  wire [63:0] _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire [511:0] _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire [63:0] _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire [511:0] _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire [63:0] _GEN_1_inputMemAddr;
  wire  _GEN_1_inputMemAddrValid;
  wire  _GEN_1_inputMemAddrReady;
  wire [511:0] _GEN_1_inputMemBlock;
  wire  _GEN_1_inputMemBlockValid;
  wire  _GEN_1_inputMemBlockReady;
  wire [63:0] _GEN_1_outputMemAddr;
  wire  _GEN_1_outputMemAddrValid;
  wire  _GEN_1_outputMemAddrReady;
  wire [511:0] _GEN_1_outputMemBlock;
  wire  _GEN_1_outputMemBlockValid;
  wire  _GEN_1_outputMemBlockReady;
  wire  _GEN_1_inputFinished;
  wire  _GEN_1_outputFinished;
  wire [63:0] _GEN_2_inputMemAddr;
  wire  _GEN_2_inputMemAddrValid;
  wire  _GEN_2_inputMemAddrReady;
  wire [511:0] _GEN_2_inputMemBlock;
  wire  _GEN_2_inputMemBlockValid;
  wire  _GEN_2_inputMemBlockReady;
  wire [63:0] _GEN_2_outputMemAddr;
  wire  _GEN_2_outputMemAddrValid;
  wire  _GEN_2_outputMemAddrReady;
  wire [511:0] _GEN_2_outputMemBlock;
  wire  _GEN_2_outputMemBlockValid;
  wire  _GEN_2_outputMemBlockReady;
  wire  _GEN_2_inputFinished;
  wire  _GEN_2_outputFinished;
  wire  _T_799;
  wire  _T_801;
  wire [511:0] _T_805;
  wire  _T_809;
  wire [63:0] _GEN_3_inputMemAddr;
  wire  _GEN_3_inputMemAddrValid;
  wire  _GEN_3_inputMemAddrReady;
  wire [511:0] _GEN_3_inputMemBlock;
  wire  _GEN_3_inputMemBlockValid;
  wire  _GEN_3_inputMemBlockReady;
  wire [63:0] _GEN_3_outputMemAddr;
  wire  _GEN_3_outputMemAddrValid;
  wire  _GEN_3_outputMemAddrReady;
  wire [511:0] _GEN_3_outputMemBlock;
  wire  _GEN_3_outputMemBlockValid;
  wire  _GEN_3_outputMemBlockReady;
  wire  _GEN_3_inputFinished;
  wire  _GEN_3_outputFinished;
  wire [63:0] _GEN_4_inputMemAddr;
  wire  _GEN_4_inputMemAddrValid;
  wire  _GEN_4_inputMemAddrReady;
  wire [511:0] _GEN_4_inputMemBlock;
  wire  _GEN_4_inputMemBlockValid;
  wire  _GEN_4_inputMemBlockReady;
  wire [63:0] _GEN_4_outputMemAddr;
  wire  _GEN_4_outputMemAddrValid;
  wire  _GEN_4_outputMemAddrReady;
  wire [511:0] _GEN_4_outputMemBlock;
  wire  _GEN_4_outputMemBlockValid;
  wire  _GEN_4_outputMemBlockReady;
  wire  _GEN_4_inputFinished;
  wire  _GEN_4_outputFinished;
  wire  _T_1068;
  wire [63:0] _GEN_5_inputMemAddr;
  wire  _GEN_5_inputMemAddrValid;
  wire  _GEN_5_inputMemAddrReady;
  wire [511:0] _GEN_5_inputMemBlock;
  wire  _GEN_5_inputMemBlockValid;
  wire  _GEN_5_inputMemBlockReady;
  wire [63:0] _GEN_5_outputMemAddr;
  wire  _GEN_5_outputMemAddrValid;
  wire  _GEN_5_outputMemAddrReady;
  wire [511:0] _GEN_5_outputMemBlock;
  wire  _GEN_5_outputMemBlockValid;
  wire  _GEN_5_outputMemBlockReady;
  wire  _GEN_5_inputFinished;
  wire  _GEN_5_outputFinished;
  wire  _T_1069;
  wire [1:0] _T_1074;
  wire  _T_1075;
  wire  _T_1076;
  wire  _GEN_54;
  wire [63:0] _GEN_6_inputMemAddr;
  wire  _GEN_6_inputMemAddrValid;
  wire  _GEN_6_inputMemAddrReady;
  wire [511:0] _GEN_6_inputMemBlock;
  wire  _GEN_6_inputMemBlockValid;
  wire  _GEN_6_inputMemBlockReady;
  wire [63:0] _GEN_6_outputMemAddr;
  wire  _GEN_6_outputMemAddrValid;
  wire  _GEN_6_outputMemAddrReady;
  wire [511:0] _GEN_6_outputMemBlock;
  wire  _GEN_6_outputMemBlockValid;
  wire  _GEN_6_outputMemBlockReady;
  wire  _GEN_6_inputFinished;
  wire  _GEN_6_outputFinished;
  wire [63:0] _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire [511:0] _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire [63:0] _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire [511:0] _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire [63:0] _GEN_7_inputMemAddr;
  wire  _GEN_7_inputMemAddrValid;
  wire  _GEN_7_inputMemAddrReady;
  wire [511:0] _GEN_7_inputMemBlock;
  wire  _GEN_7_inputMemBlockValid;
  wire  _GEN_7_inputMemBlockReady;
  wire [63:0] _GEN_7_outputMemAddr;
  wire  _GEN_7_outputMemAddrValid;
  wire  _GEN_7_outputMemAddrReady;
  wire [511:0] _GEN_7_outputMemBlock;
  wire  _GEN_7_outputMemBlockValid;
  wire  _GEN_7_outputMemBlockReady;
  wire  _GEN_7_inputFinished;
  wire  _GEN_7_outputFinished;
  wire [63:0] _GEN_8_inputMemAddr;
  wire  _GEN_8_inputMemAddrValid;
  wire  _GEN_8_inputMemAddrReady;
  wire [511:0] _GEN_8_inputMemBlock;
  wire  _GEN_8_inputMemBlockValid;
  wire  _GEN_8_inputMemBlockReady;
  wire [63:0] _GEN_8_outputMemAddr;
  wire  _GEN_8_outputMemAddrValid;
  wire  _GEN_8_outputMemAddrReady;
  wire [511:0] _GEN_8_outputMemBlock;
  wire  _GEN_8_outputMemBlockValid;
  wire  _GEN_8_outputMemBlockReady;
  wire  _GEN_8_inputFinished;
  wire  _GEN_8_outputFinished;
  wire  _T_1338;
  wire [511:0] _T_1342;
  wire  _T_1346;
  wire [63:0] _GEN_9_inputMemAddr;
  wire  _GEN_9_inputMemAddrValid;
  wire  _GEN_9_inputMemAddrReady;
  wire [511:0] _GEN_9_inputMemBlock;
  wire  _GEN_9_inputMemBlockValid;
  wire  _GEN_9_inputMemBlockReady;
  wire [63:0] _GEN_9_outputMemAddr;
  wire  _GEN_9_outputMemAddrValid;
  wire  _GEN_9_outputMemAddrReady;
  wire [511:0] _GEN_9_outputMemBlock;
  wire  _GEN_9_outputMemBlockValid;
  wire  _GEN_9_outputMemBlockReady;
  wire  _GEN_9_inputFinished;
  wire  _GEN_9_outputFinished;
  wire [63:0] _GEN_10_inputMemAddr;
  wire  _GEN_10_inputMemAddrValid;
  wire  _GEN_10_inputMemAddrReady;
  wire [511:0] _GEN_10_inputMemBlock;
  wire  _GEN_10_inputMemBlockValid;
  wire  _GEN_10_inputMemBlockReady;
  wire [63:0] _GEN_10_outputMemAddr;
  wire  _GEN_10_outputMemAddrValid;
  wire  _GEN_10_outputMemAddrReady;
  wire [511:0] _GEN_10_outputMemBlock;
  wire  _GEN_10_outputMemBlockValid;
  wire  _GEN_10_outputMemBlockReady;
  wire  _GEN_10_inputFinished;
  wire  _GEN_10_outputFinished;
  wire  _T_1605;
  wire [63:0] _GEN_11_inputMemAddr;
  wire  _GEN_11_inputMemAddrValid;
  wire  _GEN_11_inputMemAddrReady;
  wire [511:0] _GEN_11_inputMemBlock;
  wire  _GEN_11_inputMemBlockValid;
  wire  _GEN_11_inputMemBlockReady;
  wire [63:0] _GEN_11_outputMemAddr;
  wire  _GEN_11_outputMemAddrValid;
  wire  _GEN_11_outputMemAddrReady;
  wire [511:0] _GEN_11_outputMemBlock;
  wire  _GEN_11_outputMemBlockValid;
  wire  _GEN_11_outputMemBlockReady;
  wire  _GEN_11_inputFinished;
  wire  _GEN_11_outputFinished;
  wire  _T_1606;
  wire [1:0] _T_1611;
  wire  _T_1612;
  wire  _T_1613;
  wire  _GEN_83;
  wire [63:0] _GEN_12_inputMemAddr;
  wire  _GEN_12_inputMemAddrValid;
  wire  _GEN_12_inputMemAddrReady;
  wire [511:0] _GEN_12_inputMemBlock;
  wire  _GEN_12_inputMemBlockValid;
  wire  _GEN_12_inputMemBlockReady;
  wire [63:0] _GEN_12_outputMemAddr;
  wire  _GEN_12_outputMemAddrValid;
  wire  _GEN_12_outputMemAddrReady;
  wire [511:0] _GEN_12_outputMemBlock;
  wire  _GEN_12_outputMemBlockValid;
  wire  _GEN_12_outputMemBlockReady;
  wire  _GEN_12_inputFinished;
  wire  _GEN_12_outputFinished;
  wire [63:0] _GEN_84;
  wire  _GEN_85;
  wire  _GEN_86;
  wire [511:0] _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire [63:0] _GEN_90;
  wire  _GEN_91;
  wire  _GEN_92;
  wire [511:0] _GEN_93;
  wire  _GEN_94;
  wire  _GEN_95;
  wire  _GEN_96;
  wire  _GEN_97;
  wire [63:0] _GEN_13_inputMemAddr;
  wire  _GEN_13_inputMemAddrValid;
  wire  _GEN_13_inputMemAddrReady;
  wire [511:0] _GEN_13_inputMemBlock;
  wire  _GEN_13_inputMemBlockValid;
  wire  _GEN_13_inputMemBlockReady;
  wire [63:0] _GEN_13_outputMemAddr;
  wire  _GEN_13_outputMemAddrValid;
  wire  _GEN_13_outputMemAddrReady;
  wire [511:0] _GEN_13_outputMemBlock;
  wire  _GEN_13_outputMemBlockValid;
  wire  _GEN_13_outputMemBlockReady;
  wire  _GEN_13_inputFinished;
  wire  _GEN_13_outputFinished;
  wire [63:0] _GEN_14_inputMemAddr;
  wire  _GEN_14_inputMemAddrValid;
  wire  _GEN_14_inputMemAddrReady;
  wire [511:0] _GEN_14_inputMemBlock;
  wire  _GEN_14_inputMemBlockValid;
  wire  _GEN_14_inputMemBlockReady;
  wire [63:0] _GEN_14_outputMemAddr;
  wire  _GEN_14_outputMemAddrValid;
  wire  _GEN_14_outputMemAddrReady;
  wire [511:0] _GEN_14_outputMemBlock;
  wire  _GEN_14_outputMemBlockValid;
  wire  _GEN_14_outputMemBlockReady;
  wire  _GEN_14_inputFinished;
  wire  _GEN_14_outputFinished;
  wire [63:0] _GEN_15_inputMemAddr;
  wire  _GEN_15_inputMemAddrValid;
  wire  _GEN_15_inputMemAddrReady;
  wire [511:0] _GEN_15_inputMemBlock;
  wire  _GEN_15_inputMemBlockValid;
  wire  _GEN_15_inputMemBlockReady;
  wire [63:0] _GEN_15_outputMemAddr;
  wire  _GEN_15_outputMemAddrValid;
  wire  _GEN_15_outputMemAddrReady;
  wire [511:0] _GEN_15_outputMemBlock;
  wire  _GEN_15_outputMemBlockValid;
  wire  _GEN_15_outputMemBlockReady;
  wire  _GEN_15_inputFinished;
  wire  _GEN_15_outputFinished;
  wire  _T_1959;
  wire  _T_1961;
  wire  _T_1965;
  wire [63:0] _GEN_16_inputMemAddr;
  wire  _GEN_16_inputMemAddrValid;
  wire  _GEN_16_inputMemAddrReady;
  wire [511:0] _GEN_16_inputMemBlock;
  wire  _GEN_16_inputMemBlockValid;
  wire  _GEN_16_inputMemBlockReady;
  wire [63:0] _GEN_16_outputMemAddr;
  wire  _GEN_16_outputMemAddrValid;
  wire  _GEN_16_outputMemAddrReady;
  wire [511:0] _GEN_16_outputMemBlock;
  wire  _GEN_16_outputMemBlockValid;
  wire  _GEN_16_outputMemBlockReady;
  wire  _GEN_16_inputFinished;
  wire  _GEN_16_outputFinished;
  wire [63:0] _GEN_17_inputMemAddr;
  wire  _GEN_17_inputMemAddrValid;
  wire  _GEN_17_inputMemAddrReady;
  wire [511:0] _GEN_17_inputMemBlock;
  wire  _GEN_17_inputMemBlockValid;
  wire  _GEN_17_inputMemBlockReady;
  wire [63:0] _GEN_17_outputMemAddr;
  wire  _GEN_17_outputMemAddrValid;
  wire  _GEN_17_outputMemAddrReady;
  wire [511:0] _GEN_17_outputMemBlock;
  wire  _GEN_17_outputMemBlockValid;
  wire  _GEN_17_outputMemBlockReady;
  wire  _GEN_17_inputFinished;
  wire  _GEN_17_outputFinished;
  wire  _T_2224;
  wire [63:0] _GEN_18_inputMemAddr;
  wire  _GEN_18_inputMemAddrValid;
  wire  _GEN_18_inputMemAddrReady;
  wire [511:0] _GEN_18_inputMemBlock;
  wire  _GEN_18_inputMemBlockValid;
  wire  _GEN_18_inputMemBlockReady;
  wire [63:0] _GEN_18_outputMemAddr;
  wire  _GEN_18_outputMemAddrValid;
  wire  _GEN_18_outputMemAddrReady;
  wire [511:0] _GEN_18_outputMemBlock;
  wire  _GEN_18_outputMemBlockValid;
  wire  _GEN_18_outputMemBlockReady;
  wire  _GEN_18_inputFinished;
  wire  _GEN_18_outputFinished;
  wire  _T_2225;
  wire [1:0] _T_2230;
  wire  _T_2231;
  wire  _T_2232;
  wire  _GEN_112;
  wire [63:0] _GEN_19_inputMemAddr;
  wire  _GEN_19_inputMemAddrValid;
  wire  _GEN_19_inputMemAddrReady;
  wire [511:0] _GEN_19_inputMemBlock;
  wire  _GEN_19_inputMemBlockValid;
  wire  _GEN_19_inputMemBlockReady;
  wire [63:0] _GEN_19_outputMemAddr;
  wire  _GEN_19_outputMemAddrValid;
  wire  _GEN_19_outputMemAddrReady;
  wire [511:0] _GEN_19_outputMemBlock;
  wire  _GEN_19_outputMemBlockValid;
  wire  _GEN_19_outputMemBlockReady;
  wire  _GEN_19_inputFinished;
  wire  _GEN_19_outputFinished;
  wire [63:0] _GEN_113;
  wire  _GEN_114;
  wire  _GEN_115;
  wire [511:0] _GEN_116;
  wire  _GEN_117;
  wire  _GEN_118;
  wire [63:0] _GEN_119;
  wire  _GEN_120;
  wire  _GEN_121;
  wire [511:0] _GEN_122;
  wire  _GEN_123;
  wire  _GEN_124;
  wire  _GEN_125;
  wire  _GEN_126;
  wire [63:0] _GEN_20_inputMemAddr;
  wire  _GEN_20_inputMemAddrValid;
  wire  _GEN_20_inputMemAddrReady;
  wire [511:0] _GEN_20_inputMemBlock;
  wire  _GEN_20_inputMemBlockValid;
  wire  _GEN_20_inputMemBlockReady;
  wire [63:0] _GEN_20_outputMemAddr;
  wire  _GEN_20_outputMemAddrValid;
  wire  _GEN_20_outputMemAddrReady;
  wire [511:0] _GEN_20_outputMemBlock;
  wire  _GEN_20_outputMemBlockValid;
  wire  _GEN_20_outputMemBlockReady;
  wire  _GEN_20_inputFinished;
  wire  _GEN_20_outputFinished;
  wire [63:0] _GEN_21_inputMemAddr;
  wire  _GEN_21_inputMemAddrValid;
  wire  _GEN_21_inputMemAddrReady;
  wire [511:0] _GEN_21_inputMemBlock;
  wire  _GEN_21_inputMemBlockValid;
  wire  _GEN_21_inputMemBlockReady;
  wire [63:0] _GEN_21_outputMemAddr;
  wire  _GEN_21_outputMemAddrValid;
  wire  _GEN_21_outputMemAddrReady;
  wire [511:0] _GEN_21_outputMemBlock;
  wire  _GEN_21_outputMemBlockValid;
  wire  _GEN_21_outputMemBlockReady;
  wire  _GEN_21_inputFinished;
  wire  _GEN_21_outputFinished;
  wire [63:0] _GEN_22_inputMemAddr;
  wire  _GEN_22_inputMemAddrValid;
  wire  _GEN_22_inputMemAddrReady;
  wire [511:0] _GEN_22_inputMemBlock;
  wire  _GEN_22_inputMemBlockValid;
  wire  _GEN_22_inputMemBlockReady;
  wire [63:0] _GEN_22_outputMemAddr;
  wire  _GEN_22_outputMemAddrValid;
  wire  _GEN_22_outputMemAddrReady;
  wire [511:0] _GEN_22_outputMemBlock;
  wire  _GEN_22_outputMemBlockValid;
  wire  _GEN_22_outputMemBlockReady;
  wire  _GEN_22_inputFinished;
  wire  _GEN_22_outputFinished;
  wire  _T_2580;
  wire  _T_2584;
  wire [63:0] _GEN_23_inputMemAddr;
  wire  _GEN_23_inputMemAddrValid;
  wire  _GEN_23_inputMemAddrReady;
  wire [511:0] _GEN_23_inputMemBlock;
  wire  _GEN_23_inputMemBlockValid;
  wire  _GEN_23_inputMemBlockReady;
  wire [63:0] _GEN_23_outputMemAddr;
  wire  _GEN_23_outputMemAddrValid;
  wire  _GEN_23_outputMemAddrReady;
  wire [511:0] _GEN_23_outputMemBlock;
  wire  _GEN_23_outputMemBlockValid;
  wire  _GEN_23_outputMemBlockReady;
  wire  _GEN_23_inputFinished;
  wire  _GEN_23_outputFinished;
  wire [63:0] _GEN_24_inputMemAddr;
  wire  _GEN_24_inputMemAddrValid;
  wire  _GEN_24_inputMemAddrReady;
  wire [511:0] _GEN_24_inputMemBlock;
  wire  _GEN_24_inputMemBlockValid;
  wire  _GEN_24_inputMemBlockReady;
  wire [63:0] _GEN_24_outputMemAddr;
  wire  _GEN_24_outputMemAddrValid;
  wire  _GEN_24_outputMemAddrReady;
  wire [511:0] _GEN_24_outputMemBlock;
  wire  _GEN_24_outputMemBlockValid;
  wire  _GEN_24_outputMemBlockReady;
  wire  _GEN_24_inputFinished;
  wire  _GEN_24_outputFinished;
  wire  _T_2843;
  wire [63:0] _GEN_25_inputMemAddr;
  wire  _GEN_25_inputMemAddrValid;
  wire  _GEN_25_inputMemAddrReady;
  wire [511:0] _GEN_25_inputMemBlock;
  wire  _GEN_25_inputMemBlockValid;
  wire  _GEN_25_inputMemBlockReady;
  wire [63:0] _GEN_25_outputMemAddr;
  wire  _GEN_25_outputMemAddrValid;
  wire  _GEN_25_outputMemAddrReady;
  wire [511:0] _GEN_25_outputMemBlock;
  wire  _GEN_25_outputMemBlockValid;
  wire  _GEN_25_outputMemBlockReady;
  wire  _GEN_25_inputFinished;
  wire  _GEN_25_outputFinished;
  wire  _T_2844;
  wire [1:0] _T_2849;
  wire  _T_2850;
  wire  _T_2851;
  wire  _GEN_141;
  wire  cumFinished;
  StreamingCore StreamingCore (
    .clock(StreamingCore_clock),
    .reset(StreamingCore_reset),
    .io_inputMemAddr(StreamingCore_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_io_inputMemAddrValid),
    .io_inputMemAddrReady(StreamingCore_io_inputMemAddrReady),
    .io_inputMemBlock(StreamingCore_io_inputMemBlock),
    .io_inputMemBlockValid(StreamingCore_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_io_outputMemBlock),
    .io_outputMemBlockValid(StreamingCore_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_io_outputMemBlockReady),
    .io_inputFinished(StreamingCore_io_inputFinished),
    .io_outputFinished(StreamingCore_io_outputFinished)
  );
  StreamingCore_1 StreamingCore_1 (
    .clock(StreamingCore_1_clock),
    .reset(StreamingCore_1_reset),
    .io_inputMemAddr(StreamingCore_1_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_1_io_inputMemAddrValid),
    .io_inputMemAddrReady(StreamingCore_1_io_inputMemAddrReady),
    .io_inputMemBlock(StreamingCore_1_io_inputMemBlock),
    .io_inputMemBlockValid(StreamingCore_1_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_1_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_1_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_1_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_1_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_1_io_outputMemBlock),
    .io_outputMemBlockValid(StreamingCore_1_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_1_io_outputMemBlockReady),
    .io_inputFinished(StreamingCore_1_io_inputFinished),
    .io_outputFinished(StreamingCore_1_io_outputFinished)
  );
  assign io_inputMemAddrs_0 = _GEN_0_inputMemAddr;
  assign io_inputMemAddrs_1 = _GEN_6_inputMemAddr;
  assign io_inputMemAddrValids_0 = _GEN_1_inputMemAddrValid;
  assign io_inputMemAddrValids_1 = _GEN_7_inputMemAddrValid;
  assign io_inputMemBlockReadys_0 = _GEN_2_inputMemBlockReady;
  assign io_inputMemBlockReadys_1 = _GEN_8_inputMemBlockReady;
  assign io_outputMemAddrs_0 = _GEN_12_outputMemAddr;
  assign io_outputMemAddrs_1 = _GEN_19_outputMemAddr;
  assign io_outputMemAddrValids_0 = _GEN_13_outputMemAddrValid;
  assign io_outputMemAddrValids_1 = _GEN_20_outputMemAddrValid;
  assign io_outputMemBlocks_0 = _GEN_14_outputMemBlock;
  assign io_outputMemBlocks_1 = _GEN_21_outputMemBlock;
  assign io_outputMemBlockValids_0 = _GEN_15_outputMemBlockValid;
  assign io_outputMemBlockValids_1 = _GEN_22_outputMemBlockValid;
  assign io_finished = cumFinished;
  assign StreamingCore_clock = clock;
  assign StreamingCore_reset = reset;
  assign StreamingCore_io_inputMemAddrReady = cores_0_inputMemAddrReady;
  assign StreamingCore_io_inputMemBlock = cores_0_inputMemBlock;
  assign StreamingCore_io_inputMemBlockValid = cores_0_inputMemBlockValid;
  assign StreamingCore_io_outputMemAddrReady = cores_0_outputMemAddrReady;
  assign StreamingCore_io_outputMemBlockReady = cores_0_outputMemBlockReady;
  assign StreamingCore_1_clock = clock;
  assign StreamingCore_1_reset = reset;
  assign StreamingCore_1_io_inputMemAddrReady = cores_1_inputMemAddrReady;
  assign StreamingCore_1_io_inputMemBlock = cores_1_inputMemBlock;
  assign StreamingCore_1_io_inputMemBlockValid = cores_1_inputMemBlockValid;
  assign StreamingCore_1_io_outputMemAddrReady = cores_1_outputMemAddrReady;
  assign StreamingCore_1_io_outputMemBlockReady = cores_1_outputMemBlockReady;
  assign cores_0_inputMemAddr = StreamingCore_io_inputMemAddr;
  assign cores_0_inputMemAddrValid = StreamingCore_io_inputMemAddrValid;
  assign cores_0_inputMemAddrReady = _T_801;
  assign cores_0_inputMemBlock = _T_805;
  assign cores_0_inputMemBlockValid = _T_809;
  assign cores_0_inputMemBlockReady = StreamingCore_io_inputMemBlockReady;
  assign cores_0_outputMemAddr = StreamingCore_io_outputMemAddr;
  assign cores_0_outputMemAddrValid = StreamingCore_io_outputMemAddrValid;
  assign cores_0_outputMemAddrReady = _T_1961;
  assign cores_0_outputMemBlock = StreamingCore_io_outputMemBlock;
  assign cores_0_outputMemBlockValid = StreamingCore_io_outputMemBlockValid;
  assign cores_0_outputMemBlockReady = _T_1965;
  assign cores_0_inputFinished = StreamingCore_io_inputFinished;
  assign cores_0_outputFinished = StreamingCore_io_outputFinished;
  assign cores_1_inputMemAddr = StreamingCore_1_io_inputMemAddr;
  assign cores_1_inputMemAddrValid = StreamingCore_1_io_inputMemAddrValid;
  assign cores_1_inputMemAddrReady = _T_1338;
  assign cores_1_inputMemBlock = _T_1342;
  assign cores_1_inputMemBlockValid = _T_1346;
  assign cores_1_inputMemBlockReady = StreamingCore_1_io_inputMemBlockReady;
  assign cores_1_outputMemAddr = StreamingCore_1_io_outputMemAddr;
  assign cores_1_outputMemAddrValid = StreamingCore_1_io_outputMemAddrValid;
  assign cores_1_outputMemAddrReady = _T_2580;
  assign cores_1_outputMemBlock = StreamingCore_1_io_outputMemBlock;
  assign cores_1_outputMemBlockValid = StreamingCore_1_io_outputMemBlockValid;
  assign cores_1_outputMemBlockReady = _T_2584;
  assign cores_1_inputFinished = StreamingCore_1_io_inputFinished;
  assign cores_1_outputFinished = StreamingCore_1_io_outputFinished;
  assign _GEN_0_inputMemAddr = _GEN_26;
  assign _GEN_0_inputMemAddrValid = _GEN_27;
  assign _GEN_0_inputMemAddrReady = _GEN_28;
  assign _GEN_0_inputMemBlock = _GEN_29;
  assign _GEN_0_inputMemBlockValid = _GEN_30;
  assign _GEN_0_inputMemBlockReady = _GEN_31;
  assign _GEN_0_outputMemAddr = _GEN_32;
  assign _GEN_0_outputMemAddrValid = _GEN_33;
  assign _GEN_0_outputMemAddrReady = _GEN_34;
  assign _GEN_0_outputMemBlock = _GEN_35;
  assign _GEN_0_outputMemBlockValid = _GEN_36;
  assign _GEN_0_outputMemBlockReady = _GEN_37;
  assign _GEN_0_inputFinished = _GEN_38;
  assign _GEN_0_outputFinished = _GEN_39;
  assign _GEN_26 = _T_533 ? cores_1_inputMemAddr : cores_0_inputMemAddr;
  assign _GEN_27 = _T_533 ? cores_1_inputMemAddrValid : cores_0_inputMemAddrValid;
  assign _GEN_28 = _T_533 ? cores_1_inputMemAddrReady : cores_0_inputMemAddrReady;
  assign _GEN_29 = _T_533 ? cores_1_inputMemBlock : cores_0_inputMemBlock;
  assign _GEN_30 = _T_533 ? cores_1_inputMemBlockValid : cores_0_inputMemBlockValid;
  assign _GEN_31 = _T_533 ? cores_1_inputMemBlockReady : cores_0_inputMemBlockReady;
  assign _GEN_32 = _T_533 ? cores_1_outputMemAddr : cores_0_outputMemAddr;
  assign _GEN_33 = _T_533 ? cores_1_outputMemAddrValid : cores_0_outputMemAddrValid;
  assign _GEN_34 = _T_533 ? cores_1_outputMemAddrReady : cores_0_outputMemAddrReady;
  assign _GEN_35 = _T_533 ? cores_1_outputMemBlock : cores_0_outputMemBlock;
  assign _GEN_36 = _T_533 ? cores_1_outputMemBlockValid : cores_0_outputMemBlockValid;
  assign _GEN_37 = _T_533 ? cores_1_outputMemBlockReady : cores_0_outputMemBlockReady;
  assign _GEN_38 = _T_533 ? cores_1_inputFinished : cores_0_inputFinished;
  assign _GEN_39 = _T_533 ? cores_1_outputFinished : cores_0_outputFinished;
  assign _GEN_1_inputMemAddr = _GEN_26;
  assign _GEN_1_inputMemAddrValid = _GEN_27;
  assign _GEN_1_inputMemAddrReady = _GEN_28;
  assign _GEN_1_inputMemBlock = _GEN_29;
  assign _GEN_1_inputMemBlockValid = _GEN_30;
  assign _GEN_1_inputMemBlockReady = _GEN_31;
  assign _GEN_1_outputMemAddr = _GEN_32;
  assign _GEN_1_outputMemAddrValid = _GEN_33;
  assign _GEN_1_outputMemAddrReady = _GEN_34;
  assign _GEN_1_outputMemBlock = _GEN_35;
  assign _GEN_1_outputMemBlockValid = _GEN_36;
  assign _GEN_1_outputMemBlockReady = _GEN_37;
  assign _GEN_1_inputFinished = _GEN_38;
  assign _GEN_1_outputFinished = _GEN_39;
  assign _GEN_2_inputMemAddr = _GEN_26;
  assign _GEN_2_inputMemAddrValid = _GEN_27;
  assign _GEN_2_inputMemAddrReady = _GEN_28;
  assign _GEN_2_inputMemBlock = _GEN_29;
  assign _GEN_2_inputMemBlockValid = _GEN_30;
  assign _GEN_2_inputMemBlockReady = _GEN_31;
  assign _GEN_2_outputMemAddr = _GEN_32;
  assign _GEN_2_outputMemAddrValid = _GEN_33;
  assign _GEN_2_outputMemAddrReady = _GEN_34;
  assign _GEN_2_outputMemBlock = _GEN_35;
  assign _GEN_2_outputMemBlockValid = _GEN_36;
  assign _GEN_2_outputMemBlockReady = _GEN_37;
  assign _GEN_2_inputFinished = _GEN_38;
  assign _GEN_2_outputFinished = _GEN_39;
  assign _T_799 = _T_533 == 1'h0;
  assign _T_801 = _T_799 ? io_inputMemAddrReadys_0 : 1'h0;
  assign _T_805 = _T_799 ? io_inputMemBlocks_0 : 512'h0;
  assign _T_809 = _T_799 ? io_inputMemBlockValids_0 : 1'h0;
  assign _GEN_3_inputMemAddr = _GEN_26;
  assign _GEN_3_inputMemAddrValid = _GEN_27;
  assign _GEN_3_inputMemAddrReady = _GEN_28;
  assign _GEN_3_inputMemBlock = _GEN_29;
  assign _GEN_3_inputMemBlockValid = _GEN_30;
  assign _GEN_3_inputMemBlockReady = _GEN_31;
  assign _GEN_3_outputMemAddr = _GEN_32;
  assign _GEN_3_outputMemAddrValid = _GEN_33;
  assign _GEN_3_outputMemAddrReady = _GEN_34;
  assign _GEN_3_outputMemBlock = _GEN_35;
  assign _GEN_3_outputMemBlockValid = _GEN_36;
  assign _GEN_3_outputMemBlockReady = _GEN_37;
  assign _GEN_3_inputFinished = _GEN_38;
  assign _GEN_3_outputFinished = _GEN_39;
  assign _GEN_4_inputMemAddr = _GEN_26;
  assign _GEN_4_inputMemAddrValid = _GEN_27;
  assign _GEN_4_inputMemAddrReady = _GEN_28;
  assign _GEN_4_inputMemBlock = _GEN_29;
  assign _GEN_4_inputMemBlockValid = _GEN_30;
  assign _GEN_4_inputMemBlockReady = _GEN_31;
  assign _GEN_4_outputMemAddr = _GEN_32;
  assign _GEN_4_outputMemAddrValid = _GEN_33;
  assign _GEN_4_outputMemAddrReady = _GEN_34;
  assign _GEN_4_outputMemBlock = _GEN_35;
  assign _GEN_4_outputMemBlockValid = _GEN_36;
  assign _GEN_4_outputMemBlockReady = _GEN_37;
  assign _GEN_4_inputFinished = _GEN_38;
  assign _GEN_4_outputFinished = _GEN_39;
  assign _T_1068 = _GEN_3_inputMemBlockReady & _GEN_4_inputMemBlockValid;
  assign _GEN_5_inputMemAddr = _GEN_26;
  assign _GEN_5_inputMemAddrValid = _GEN_27;
  assign _GEN_5_inputMemAddrReady = _GEN_28;
  assign _GEN_5_inputMemBlock = _GEN_29;
  assign _GEN_5_inputMemBlockValid = _GEN_30;
  assign _GEN_5_inputMemBlockReady = _GEN_31;
  assign _GEN_5_outputMemAddr = _GEN_32;
  assign _GEN_5_outputMemAddrValid = _GEN_33;
  assign _GEN_5_outputMemAddrReady = _GEN_34;
  assign _GEN_5_outputMemBlock = _GEN_35;
  assign _GEN_5_outputMemBlockValid = _GEN_36;
  assign _GEN_5_outputMemBlockReady = _GEN_37;
  assign _GEN_5_inputFinished = _GEN_38;
  assign _GEN_5_outputFinished = _GEN_39;
  assign _T_1069 = _GEN_5_inputFinished | _T_1068;
  assign _T_1074 = _T_533 + 1'h1;
  assign _T_1075 = _T_1074[0:0];
  assign _T_1076 = _T_799 ? 1'h0 : _T_1075;
  assign _GEN_54 = _T_1069 ? _T_1076 : _T_533;
  assign _GEN_6_inputMemAddr = _GEN_55;
  assign _GEN_6_inputMemAddrValid = _GEN_56;
  assign _GEN_6_inputMemAddrReady = _GEN_57;
  assign _GEN_6_inputMemBlock = _GEN_58;
  assign _GEN_6_inputMemBlockValid = _GEN_59;
  assign _GEN_6_inputMemBlockReady = _GEN_60;
  assign _GEN_6_outputMemAddr = _GEN_61;
  assign _GEN_6_outputMemAddrValid = _GEN_62;
  assign _GEN_6_outputMemAddrReady = _GEN_63;
  assign _GEN_6_outputMemBlock = _GEN_64;
  assign _GEN_6_outputMemBlockValid = _GEN_65;
  assign _GEN_6_outputMemBlockReady = _GEN_66;
  assign _GEN_6_inputFinished = _GEN_67;
  assign _GEN_6_outputFinished = _GEN_68;
  assign _GEN_55 = _T_535 ? cores_1_inputMemAddr : cores_0_inputMemAddr;
  assign _GEN_56 = _T_535 ? cores_1_inputMemAddrValid : cores_0_inputMemAddrValid;
  assign _GEN_57 = _T_535 ? cores_1_inputMemAddrReady : cores_0_inputMemAddrReady;
  assign _GEN_58 = _T_535 ? cores_1_inputMemBlock : cores_0_inputMemBlock;
  assign _GEN_59 = _T_535 ? cores_1_inputMemBlockValid : cores_0_inputMemBlockValid;
  assign _GEN_60 = _T_535 ? cores_1_inputMemBlockReady : cores_0_inputMemBlockReady;
  assign _GEN_61 = _T_535 ? cores_1_outputMemAddr : cores_0_outputMemAddr;
  assign _GEN_62 = _T_535 ? cores_1_outputMemAddrValid : cores_0_outputMemAddrValid;
  assign _GEN_63 = _T_535 ? cores_1_outputMemAddrReady : cores_0_outputMemAddrReady;
  assign _GEN_64 = _T_535 ? cores_1_outputMemBlock : cores_0_outputMemBlock;
  assign _GEN_65 = _T_535 ? cores_1_outputMemBlockValid : cores_0_outputMemBlockValid;
  assign _GEN_66 = _T_535 ? cores_1_outputMemBlockReady : cores_0_outputMemBlockReady;
  assign _GEN_67 = _T_535 ? cores_1_inputFinished : cores_0_inputFinished;
  assign _GEN_68 = _T_535 ? cores_1_outputFinished : cores_0_outputFinished;
  assign _GEN_7_inputMemAddr = _GEN_55;
  assign _GEN_7_inputMemAddrValid = _GEN_56;
  assign _GEN_7_inputMemAddrReady = _GEN_57;
  assign _GEN_7_inputMemBlock = _GEN_58;
  assign _GEN_7_inputMemBlockValid = _GEN_59;
  assign _GEN_7_inputMemBlockReady = _GEN_60;
  assign _GEN_7_outputMemAddr = _GEN_61;
  assign _GEN_7_outputMemAddrValid = _GEN_62;
  assign _GEN_7_outputMemAddrReady = _GEN_63;
  assign _GEN_7_outputMemBlock = _GEN_64;
  assign _GEN_7_outputMemBlockValid = _GEN_65;
  assign _GEN_7_outputMemBlockReady = _GEN_66;
  assign _GEN_7_inputFinished = _GEN_67;
  assign _GEN_7_outputFinished = _GEN_68;
  assign _GEN_8_inputMemAddr = _GEN_55;
  assign _GEN_8_inputMemAddrValid = _GEN_56;
  assign _GEN_8_inputMemAddrReady = _GEN_57;
  assign _GEN_8_inputMemBlock = _GEN_58;
  assign _GEN_8_inputMemBlockValid = _GEN_59;
  assign _GEN_8_inputMemBlockReady = _GEN_60;
  assign _GEN_8_outputMemAddr = _GEN_61;
  assign _GEN_8_outputMemAddrValid = _GEN_62;
  assign _GEN_8_outputMemAddrReady = _GEN_63;
  assign _GEN_8_outputMemBlock = _GEN_64;
  assign _GEN_8_outputMemBlockValid = _GEN_65;
  assign _GEN_8_outputMemBlockReady = _GEN_66;
  assign _GEN_8_inputFinished = _GEN_67;
  assign _GEN_8_outputFinished = _GEN_68;
  assign _T_1338 = _T_535 ? io_inputMemAddrReadys_1 : 1'h0;
  assign _T_1342 = _T_535 ? io_inputMemBlocks_1 : 512'h0;
  assign _T_1346 = _T_535 ? io_inputMemBlockValids_1 : 1'h0;
  assign _GEN_9_inputMemAddr = _GEN_55;
  assign _GEN_9_inputMemAddrValid = _GEN_56;
  assign _GEN_9_inputMemAddrReady = _GEN_57;
  assign _GEN_9_inputMemBlock = _GEN_58;
  assign _GEN_9_inputMemBlockValid = _GEN_59;
  assign _GEN_9_inputMemBlockReady = _GEN_60;
  assign _GEN_9_outputMemAddr = _GEN_61;
  assign _GEN_9_outputMemAddrValid = _GEN_62;
  assign _GEN_9_outputMemAddrReady = _GEN_63;
  assign _GEN_9_outputMemBlock = _GEN_64;
  assign _GEN_9_outputMemBlockValid = _GEN_65;
  assign _GEN_9_outputMemBlockReady = _GEN_66;
  assign _GEN_9_inputFinished = _GEN_67;
  assign _GEN_9_outputFinished = _GEN_68;
  assign _GEN_10_inputMemAddr = _GEN_55;
  assign _GEN_10_inputMemAddrValid = _GEN_56;
  assign _GEN_10_inputMemAddrReady = _GEN_57;
  assign _GEN_10_inputMemBlock = _GEN_58;
  assign _GEN_10_inputMemBlockValid = _GEN_59;
  assign _GEN_10_inputMemBlockReady = _GEN_60;
  assign _GEN_10_outputMemAddr = _GEN_61;
  assign _GEN_10_outputMemAddrValid = _GEN_62;
  assign _GEN_10_outputMemAddrReady = _GEN_63;
  assign _GEN_10_outputMemBlock = _GEN_64;
  assign _GEN_10_outputMemBlockValid = _GEN_65;
  assign _GEN_10_outputMemBlockReady = _GEN_66;
  assign _GEN_10_inputFinished = _GEN_67;
  assign _GEN_10_outputFinished = _GEN_68;
  assign _T_1605 = _GEN_9_inputMemBlockReady & _GEN_10_inputMemBlockValid;
  assign _GEN_11_inputMemAddr = _GEN_55;
  assign _GEN_11_inputMemAddrValid = _GEN_56;
  assign _GEN_11_inputMemAddrReady = _GEN_57;
  assign _GEN_11_inputMemBlock = _GEN_58;
  assign _GEN_11_inputMemBlockValid = _GEN_59;
  assign _GEN_11_inputMemBlockReady = _GEN_60;
  assign _GEN_11_outputMemAddr = _GEN_61;
  assign _GEN_11_outputMemAddrValid = _GEN_62;
  assign _GEN_11_outputMemAddrReady = _GEN_63;
  assign _GEN_11_outputMemBlock = _GEN_64;
  assign _GEN_11_outputMemBlockValid = _GEN_65;
  assign _GEN_11_outputMemBlockReady = _GEN_66;
  assign _GEN_11_inputFinished = _GEN_67;
  assign _GEN_11_outputFinished = _GEN_68;
  assign _T_1606 = _GEN_11_inputFinished | _T_1605;
  assign _T_1611 = _T_535 + 1'h1;
  assign _T_1612 = _T_1611[0:0];
  assign _T_1613 = _T_535 ? 1'h1 : _T_1612;
  assign _GEN_83 = _T_1606 ? _T_1613 : _T_535;
  assign _GEN_12_inputMemAddr = _GEN_84;
  assign _GEN_12_inputMemAddrValid = _GEN_85;
  assign _GEN_12_inputMemAddrReady = _GEN_86;
  assign _GEN_12_inputMemBlock = _GEN_87;
  assign _GEN_12_inputMemBlockValid = _GEN_88;
  assign _GEN_12_inputMemBlockReady = _GEN_89;
  assign _GEN_12_outputMemAddr = _GEN_90;
  assign _GEN_12_outputMemAddrValid = _GEN_91;
  assign _GEN_12_outputMemAddrReady = _GEN_92;
  assign _GEN_12_outputMemBlock = _GEN_93;
  assign _GEN_12_outputMemBlockValid = _GEN_94;
  assign _GEN_12_outputMemBlockReady = _GEN_95;
  assign _GEN_12_inputFinished = _GEN_96;
  assign _GEN_12_outputFinished = _GEN_97;
  assign _GEN_84 = _T_537 ? cores_1_inputMemAddr : cores_0_inputMemAddr;
  assign _GEN_85 = _T_537 ? cores_1_inputMemAddrValid : cores_0_inputMemAddrValid;
  assign _GEN_86 = _T_537 ? cores_1_inputMemAddrReady : cores_0_inputMemAddrReady;
  assign _GEN_87 = _T_537 ? cores_1_inputMemBlock : cores_0_inputMemBlock;
  assign _GEN_88 = _T_537 ? cores_1_inputMemBlockValid : cores_0_inputMemBlockValid;
  assign _GEN_89 = _T_537 ? cores_1_inputMemBlockReady : cores_0_inputMemBlockReady;
  assign _GEN_90 = _T_537 ? cores_1_outputMemAddr : cores_0_outputMemAddr;
  assign _GEN_91 = _T_537 ? cores_1_outputMemAddrValid : cores_0_outputMemAddrValid;
  assign _GEN_92 = _T_537 ? cores_1_outputMemAddrReady : cores_0_outputMemAddrReady;
  assign _GEN_93 = _T_537 ? cores_1_outputMemBlock : cores_0_outputMemBlock;
  assign _GEN_94 = _T_537 ? cores_1_outputMemBlockValid : cores_0_outputMemBlockValid;
  assign _GEN_95 = _T_537 ? cores_1_outputMemBlockReady : cores_0_outputMemBlockReady;
  assign _GEN_96 = _T_537 ? cores_1_inputFinished : cores_0_inputFinished;
  assign _GEN_97 = _T_537 ? cores_1_outputFinished : cores_0_outputFinished;
  assign _GEN_13_inputMemAddr = _GEN_84;
  assign _GEN_13_inputMemAddrValid = _GEN_85;
  assign _GEN_13_inputMemAddrReady = _GEN_86;
  assign _GEN_13_inputMemBlock = _GEN_87;
  assign _GEN_13_inputMemBlockValid = _GEN_88;
  assign _GEN_13_inputMemBlockReady = _GEN_89;
  assign _GEN_13_outputMemAddr = _GEN_90;
  assign _GEN_13_outputMemAddrValid = _GEN_91;
  assign _GEN_13_outputMemAddrReady = _GEN_92;
  assign _GEN_13_outputMemBlock = _GEN_93;
  assign _GEN_13_outputMemBlockValid = _GEN_94;
  assign _GEN_13_outputMemBlockReady = _GEN_95;
  assign _GEN_13_inputFinished = _GEN_96;
  assign _GEN_13_outputFinished = _GEN_97;
  assign _GEN_14_inputMemAddr = _GEN_84;
  assign _GEN_14_inputMemAddrValid = _GEN_85;
  assign _GEN_14_inputMemAddrReady = _GEN_86;
  assign _GEN_14_inputMemBlock = _GEN_87;
  assign _GEN_14_inputMemBlockValid = _GEN_88;
  assign _GEN_14_inputMemBlockReady = _GEN_89;
  assign _GEN_14_outputMemAddr = _GEN_90;
  assign _GEN_14_outputMemAddrValid = _GEN_91;
  assign _GEN_14_outputMemAddrReady = _GEN_92;
  assign _GEN_14_outputMemBlock = _GEN_93;
  assign _GEN_14_outputMemBlockValid = _GEN_94;
  assign _GEN_14_outputMemBlockReady = _GEN_95;
  assign _GEN_14_inputFinished = _GEN_96;
  assign _GEN_14_outputFinished = _GEN_97;
  assign _GEN_15_inputMemAddr = _GEN_84;
  assign _GEN_15_inputMemAddrValid = _GEN_85;
  assign _GEN_15_inputMemAddrReady = _GEN_86;
  assign _GEN_15_inputMemBlock = _GEN_87;
  assign _GEN_15_inputMemBlockValid = _GEN_88;
  assign _GEN_15_inputMemBlockReady = _GEN_89;
  assign _GEN_15_outputMemAddr = _GEN_90;
  assign _GEN_15_outputMemAddrValid = _GEN_91;
  assign _GEN_15_outputMemAddrReady = _GEN_92;
  assign _GEN_15_outputMemBlock = _GEN_93;
  assign _GEN_15_outputMemBlockValid = _GEN_94;
  assign _GEN_15_outputMemBlockReady = _GEN_95;
  assign _GEN_15_inputFinished = _GEN_96;
  assign _GEN_15_outputFinished = _GEN_97;
  assign _T_1959 = _T_537 == 1'h0;
  assign _T_1961 = _T_1959 ? io_outputMemAddrReadys_0 : 1'h0;
  assign _T_1965 = _T_1959 ? io_outputMemBlockReadys_0 : 1'h0;
  assign _GEN_16_inputMemAddr = _GEN_84;
  assign _GEN_16_inputMemAddrValid = _GEN_85;
  assign _GEN_16_inputMemAddrReady = _GEN_86;
  assign _GEN_16_inputMemBlock = _GEN_87;
  assign _GEN_16_inputMemBlockValid = _GEN_88;
  assign _GEN_16_inputMemBlockReady = _GEN_89;
  assign _GEN_16_outputMemAddr = _GEN_90;
  assign _GEN_16_outputMemAddrValid = _GEN_91;
  assign _GEN_16_outputMemAddrReady = _GEN_92;
  assign _GEN_16_outputMemBlock = _GEN_93;
  assign _GEN_16_outputMemBlockValid = _GEN_94;
  assign _GEN_16_outputMemBlockReady = _GEN_95;
  assign _GEN_16_inputFinished = _GEN_96;
  assign _GEN_16_outputFinished = _GEN_97;
  assign _GEN_17_inputMemAddr = _GEN_84;
  assign _GEN_17_inputMemAddrValid = _GEN_85;
  assign _GEN_17_inputMemAddrReady = _GEN_86;
  assign _GEN_17_inputMemBlock = _GEN_87;
  assign _GEN_17_inputMemBlockValid = _GEN_88;
  assign _GEN_17_inputMemBlockReady = _GEN_89;
  assign _GEN_17_outputMemAddr = _GEN_90;
  assign _GEN_17_outputMemAddrValid = _GEN_91;
  assign _GEN_17_outputMemAddrReady = _GEN_92;
  assign _GEN_17_outputMemBlock = _GEN_93;
  assign _GEN_17_outputMemBlockValid = _GEN_94;
  assign _GEN_17_outputMemBlockReady = _GEN_95;
  assign _GEN_17_inputFinished = _GEN_96;
  assign _GEN_17_outputFinished = _GEN_97;
  assign _T_2224 = _GEN_16_outputMemBlockReady & _GEN_17_outputMemBlockValid;
  assign _GEN_18_inputMemAddr = _GEN_84;
  assign _GEN_18_inputMemAddrValid = _GEN_85;
  assign _GEN_18_inputMemAddrReady = _GEN_86;
  assign _GEN_18_inputMemBlock = _GEN_87;
  assign _GEN_18_inputMemBlockValid = _GEN_88;
  assign _GEN_18_inputMemBlockReady = _GEN_89;
  assign _GEN_18_outputMemAddr = _GEN_90;
  assign _GEN_18_outputMemAddrValid = _GEN_91;
  assign _GEN_18_outputMemAddrReady = _GEN_92;
  assign _GEN_18_outputMemBlock = _GEN_93;
  assign _GEN_18_outputMemBlockValid = _GEN_94;
  assign _GEN_18_outputMemBlockReady = _GEN_95;
  assign _GEN_18_inputFinished = _GEN_96;
  assign _GEN_18_outputFinished = _GEN_97;
  assign _T_2225 = _GEN_18_outputFinished | _T_2224;
  assign _T_2230 = _T_537 + 1'h1;
  assign _T_2231 = _T_2230[0:0];
  assign _T_2232 = _T_1959 ? 1'h0 : _T_2231;
  assign _GEN_112 = _T_2225 ? _T_2232 : _T_537;
  assign _GEN_19_inputMemAddr = _GEN_113;
  assign _GEN_19_inputMemAddrValid = _GEN_114;
  assign _GEN_19_inputMemAddrReady = _GEN_115;
  assign _GEN_19_inputMemBlock = _GEN_116;
  assign _GEN_19_inputMemBlockValid = _GEN_117;
  assign _GEN_19_inputMemBlockReady = _GEN_118;
  assign _GEN_19_outputMemAddr = _GEN_119;
  assign _GEN_19_outputMemAddrValid = _GEN_120;
  assign _GEN_19_outputMemAddrReady = _GEN_121;
  assign _GEN_19_outputMemBlock = _GEN_122;
  assign _GEN_19_outputMemBlockValid = _GEN_123;
  assign _GEN_19_outputMemBlockReady = _GEN_124;
  assign _GEN_19_inputFinished = _GEN_125;
  assign _GEN_19_outputFinished = _GEN_126;
  assign _GEN_113 = _T_539 ? cores_1_inputMemAddr : cores_0_inputMemAddr;
  assign _GEN_114 = _T_539 ? cores_1_inputMemAddrValid : cores_0_inputMemAddrValid;
  assign _GEN_115 = _T_539 ? cores_1_inputMemAddrReady : cores_0_inputMemAddrReady;
  assign _GEN_116 = _T_539 ? cores_1_inputMemBlock : cores_0_inputMemBlock;
  assign _GEN_117 = _T_539 ? cores_1_inputMemBlockValid : cores_0_inputMemBlockValid;
  assign _GEN_118 = _T_539 ? cores_1_inputMemBlockReady : cores_0_inputMemBlockReady;
  assign _GEN_119 = _T_539 ? cores_1_outputMemAddr : cores_0_outputMemAddr;
  assign _GEN_120 = _T_539 ? cores_1_outputMemAddrValid : cores_0_outputMemAddrValid;
  assign _GEN_121 = _T_539 ? cores_1_outputMemAddrReady : cores_0_outputMemAddrReady;
  assign _GEN_122 = _T_539 ? cores_1_outputMemBlock : cores_0_outputMemBlock;
  assign _GEN_123 = _T_539 ? cores_1_outputMemBlockValid : cores_0_outputMemBlockValid;
  assign _GEN_124 = _T_539 ? cores_1_outputMemBlockReady : cores_0_outputMemBlockReady;
  assign _GEN_125 = _T_539 ? cores_1_inputFinished : cores_0_inputFinished;
  assign _GEN_126 = _T_539 ? cores_1_outputFinished : cores_0_outputFinished;
  assign _GEN_20_inputMemAddr = _GEN_113;
  assign _GEN_20_inputMemAddrValid = _GEN_114;
  assign _GEN_20_inputMemAddrReady = _GEN_115;
  assign _GEN_20_inputMemBlock = _GEN_116;
  assign _GEN_20_inputMemBlockValid = _GEN_117;
  assign _GEN_20_inputMemBlockReady = _GEN_118;
  assign _GEN_20_outputMemAddr = _GEN_119;
  assign _GEN_20_outputMemAddrValid = _GEN_120;
  assign _GEN_20_outputMemAddrReady = _GEN_121;
  assign _GEN_20_outputMemBlock = _GEN_122;
  assign _GEN_20_outputMemBlockValid = _GEN_123;
  assign _GEN_20_outputMemBlockReady = _GEN_124;
  assign _GEN_20_inputFinished = _GEN_125;
  assign _GEN_20_outputFinished = _GEN_126;
  assign _GEN_21_inputMemAddr = _GEN_113;
  assign _GEN_21_inputMemAddrValid = _GEN_114;
  assign _GEN_21_inputMemAddrReady = _GEN_115;
  assign _GEN_21_inputMemBlock = _GEN_116;
  assign _GEN_21_inputMemBlockValid = _GEN_117;
  assign _GEN_21_inputMemBlockReady = _GEN_118;
  assign _GEN_21_outputMemAddr = _GEN_119;
  assign _GEN_21_outputMemAddrValid = _GEN_120;
  assign _GEN_21_outputMemAddrReady = _GEN_121;
  assign _GEN_21_outputMemBlock = _GEN_122;
  assign _GEN_21_outputMemBlockValid = _GEN_123;
  assign _GEN_21_outputMemBlockReady = _GEN_124;
  assign _GEN_21_inputFinished = _GEN_125;
  assign _GEN_21_outputFinished = _GEN_126;
  assign _GEN_22_inputMemAddr = _GEN_113;
  assign _GEN_22_inputMemAddrValid = _GEN_114;
  assign _GEN_22_inputMemAddrReady = _GEN_115;
  assign _GEN_22_inputMemBlock = _GEN_116;
  assign _GEN_22_inputMemBlockValid = _GEN_117;
  assign _GEN_22_inputMemBlockReady = _GEN_118;
  assign _GEN_22_outputMemAddr = _GEN_119;
  assign _GEN_22_outputMemAddrValid = _GEN_120;
  assign _GEN_22_outputMemAddrReady = _GEN_121;
  assign _GEN_22_outputMemBlock = _GEN_122;
  assign _GEN_22_outputMemBlockValid = _GEN_123;
  assign _GEN_22_outputMemBlockReady = _GEN_124;
  assign _GEN_22_inputFinished = _GEN_125;
  assign _GEN_22_outputFinished = _GEN_126;
  assign _T_2580 = _T_539 ? io_outputMemAddrReadys_1 : 1'h0;
  assign _T_2584 = _T_539 ? io_outputMemBlockReadys_1 : 1'h0;
  assign _GEN_23_inputMemAddr = _GEN_113;
  assign _GEN_23_inputMemAddrValid = _GEN_114;
  assign _GEN_23_inputMemAddrReady = _GEN_115;
  assign _GEN_23_inputMemBlock = _GEN_116;
  assign _GEN_23_inputMemBlockValid = _GEN_117;
  assign _GEN_23_inputMemBlockReady = _GEN_118;
  assign _GEN_23_outputMemAddr = _GEN_119;
  assign _GEN_23_outputMemAddrValid = _GEN_120;
  assign _GEN_23_outputMemAddrReady = _GEN_121;
  assign _GEN_23_outputMemBlock = _GEN_122;
  assign _GEN_23_outputMemBlockValid = _GEN_123;
  assign _GEN_23_outputMemBlockReady = _GEN_124;
  assign _GEN_23_inputFinished = _GEN_125;
  assign _GEN_23_outputFinished = _GEN_126;
  assign _GEN_24_inputMemAddr = _GEN_113;
  assign _GEN_24_inputMemAddrValid = _GEN_114;
  assign _GEN_24_inputMemAddrReady = _GEN_115;
  assign _GEN_24_inputMemBlock = _GEN_116;
  assign _GEN_24_inputMemBlockValid = _GEN_117;
  assign _GEN_24_inputMemBlockReady = _GEN_118;
  assign _GEN_24_outputMemAddr = _GEN_119;
  assign _GEN_24_outputMemAddrValid = _GEN_120;
  assign _GEN_24_outputMemAddrReady = _GEN_121;
  assign _GEN_24_outputMemBlock = _GEN_122;
  assign _GEN_24_outputMemBlockValid = _GEN_123;
  assign _GEN_24_outputMemBlockReady = _GEN_124;
  assign _GEN_24_inputFinished = _GEN_125;
  assign _GEN_24_outputFinished = _GEN_126;
  assign _T_2843 = _GEN_23_outputMemBlockReady & _GEN_24_outputMemBlockValid;
  assign _GEN_25_inputMemAddr = _GEN_113;
  assign _GEN_25_inputMemAddrValid = _GEN_114;
  assign _GEN_25_inputMemAddrReady = _GEN_115;
  assign _GEN_25_inputMemBlock = _GEN_116;
  assign _GEN_25_inputMemBlockValid = _GEN_117;
  assign _GEN_25_inputMemBlockReady = _GEN_118;
  assign _GEN_25_outputMemAddr = _GEN_119;
  assign _GEN_25_outputMemAddrValid = _GEN_120;
  assign _GEN_25_outputMemAddrReady = _GEN_121;
  assign _GEN_25_outputMemBlock = _GEN_122;
  assign _GEN_25_outputMemBlockValid = _GEN_123;
  assign _GEN_25_outputMemBlockReady = _GEN_124;
  assign _GEN_25_inputFinished = _GEN_125;
  assign _GEN_25_outputFinished = _GEN_126;
  assign _T_2844 = _GEN_25_outputFinished | _T_2843;
  assign _T_2849 = _T_539 + 1'h1;
  assign _T_2850 = _T_2849[0:0];
  assign _T_2851 = _T_539 ? 1'h1 : _T_2850;
  assign _GEN_141 = _T_2844 ? _T_2851 : _T_539;
  assign cumFinished = cores_0_outputFinished & cores_1_outputFinished;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_0 = {1{$random}};
  _T_533 = _GEN_0[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1 = {1{$random}};
  _T_535 = _GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2 = {1{$random}};
  _T_537 = _GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_3 = {1{$random}};
  _T_539 = _GEN_3[0:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      _T_533 <= 1'h0;
    end else begin
      if (_T_1069) begin
        if (_T_799) begin
          _T_533 <= 1'h0;
        end else begin
          _T_533 <= _T_1075;
        end
      end
    end
    if (reset) begin
      _T_535 <= 1'h1;
    end else begin
      if (_T_1606) begin
        if (_T_535) begin
          _T_535 <= 1'h1;
        end else begin
          _T_535 <= _T_1612;
        end
      end
    end
    if (reset) begin
      _T_537 <= 1'h0;
    end else begin
      if (_T_2225) begin
        if (_T_1959) begin
          _T_537 <= 1'h0;
        end else begin
          _T_537 <= _T_2231;
        end
      end
    end
    if (reset) begin
      _T_539 <= 1'h1;
    end else begin
      if (_T_2844) begin
        if (_T_539) begin
          _T_539 <= 1'h1;
        end else begin
          _T_539 <= _T_2850;
        end
      end
    end
  end
endmodule
