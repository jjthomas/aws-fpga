`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module DualPortBRAM(
  input         clock,
  input  [4:0]  io_a_addr,
  input  [15:0] io_a_din,
  input         io_a_wr,
  input  [4:0]  io_b_addr,
  output [15:0] io_b_dout
);
  reg [15:0] mem [0:31];
  reg [31:0] _RAND_0;
  wire [15:0] mem__T_12_data;
  wire [4:0] mem__T_12_addr;
  wire [15:0] mem__T_14_data;
  wire [4:0] mem__T_14_addr;
  wire [15:0] mem__T_13_data;
  wire [4:0] mem__T_13_addr;
  wire  mem__T_13_mask;
  wire  mem__T_13_en;
  wire [15:0] mem__T_15_data;
  wire [4:0] mem__T_15_addr;
  wire  mem__T_15_mask;
  wire  mem__T_15_en;
  wire  _GEN_8;
  reg [4:0] mem__T_12_addr_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] mem__T_14_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign mem__T_12_addr = mem__T_12_addr_pipe_0;
  assign mem__T_12_data = mem[mem__T_12_addr];
  assign mem__T_14_addr = mem__T_14_addr_pipe_0;
  assign mem__T_14_data = mem[mem__T_14_addr];
  assign mem__T_13_data = io_a_din;
  assign mem__T_13_addr = io_a_addr;
  assign mem__T_13_mask = io_a_wr;
  assign mem__T_13_en = io_a_wr;
  assign mem__T_15_data = 16'h0;
  assign mem__T_15_addr = io_b_addr;
  assign mem__T_15_mask = 1'h0;
  assign mem__T_15_en = 1'h0;
  assign _GEN_8 = 1'h1;
  assign io_b_dout = mem__T_14_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem__T_12_addr_pipe_0 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem__T_14_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_13_en & mem__T_13_mask) begin
      mem[mem__T_13_addr] <= mem__T_13_data;
    end
    if(mem__T_15_en & mem__T_15_mask) begin
      mem[mem__T_15_addr] <= mem__T_15_data;
    end
    if (_GEN_8) begin
      mem__T_12_addr_pipe_0 <= io_a_addr;
    end
    if (_GEN_8) begin
      mem__T_14_addr_pipe_0 <= io_b_addr;
    end
  end
endmodule
module PassThrough(
  input         clock,
  input         reset,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  input  [9:0]  io_inputBits,
  output        io_inputMemConsumed,
  input         io_inputFinished,
  output [15:0] io_outputMemBlock,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output [9:0]  io_outputBits,
  output        io_outputFinished,
  input         io_outputMemFlushed
);
  reg  inputMemBlock_0;
  reg [31:0] _RAND_0;
  reg  inputMemBlock_1;
  reg [31:0] _RAND_1;
  reg  inputMemBlock_2;
  reg [31:0] _RAND_2;
  reg  inputMemBlock_3;
  reg [31:0] _RAND_3;
  reg  inputMemBlock_4;
  reg [31:0] _RAND_4;
  reg  inputMemBlock_5;
  reg [31:0] _RAND_5;
  reg  inputMemBlock_6;
  reg [31:0] _RAND_6;
  reg  inputMemBlock_7;
  reg [31:0] _RAND_7;
  reg  inputMemBlock_8;
  reg [31:0] _RAND_8;
  reg  inputMemBlock_9;
  reg [31:0] _RAND_9;
  reg  inputMemBlock_10;
  reg [31:0] _RAND_10;
  reg  inputMemBlock_11;
  reg [31:0] _RAND_11;
  reg  inputMemBlock_12;
  reg [31:0] _RAND_12;
  reg  inputMemBlock_13;
  reg [31:0] _RAND_13;
  reg  inputMemBlock_14;
  reg [31:0] _RAND_14;
  reg  inputMemBlock_15;
  reg [31:0] _RAND_15;
  reg [4:0] inputPieceBitsRemaining;
  reg [31:0] _RAND_16;
  reg [9:0] inputBitsRemaining;
  reg [31:0] _RAND_17;
  reg  inputBlockLoaded;
  reg [31:0] _RAND_18;
  reg  outputMemBlock_0;
  reg [31:0] _RAND_19;
  reg  outputMemBlock_1;
  reg [31:0] _RAND_20;
  reg  outputMemBlock_2;
  reg [31:0] _RAND_21;
  reg  outputMemBlock_3;
  reg [31:0] _RAND_22;
  reg  outputMemBlock_4;
  reg [31:0] _RAND_23;
  reg  outputMemBlock_5;
  reg [31:0] _RAND_24;
  reg  outputMemBlock_6;
  reg [31:0] _RAND_25;
  reg  outputMemBlock_7;
  reg [31:0] _RAND_26;
  reg  outputMemBlock_8;
  reg [31:0] _RAND_27;
  reg  outputMemBlock_9;
  reg [31:0] _RAND_28;
  reg  outputMemBlock_10;
  reg [31:0] _RAND_29;
  reg  outputMemBlock_11;
  reg [31:0] _RAND_30;
  reg  outputMemBlock_12;
  reg [31:0] _RAND_31;
  reg  outputMemBlock_13;
  reg [31:0] _RAND_32;
  reg  outputMemBlock_14;
  reg [31:0] _RAND_33;
  reg  outputMemBlock_15;
  reg [31:0] _RAND_34;
  reg [9:0] outputBits;
  reg [31:0] _RAND_35;
  reg [4:0] outputPieceBits;
  reg [31:0] _RAND_36;
  wire  inputBram_clock;
  wire [4:0] inputBram_io_a_addr;
  wire [15:0] inputBram_io_a_din;
  wire  inputBram_io_a_wr;
  wire [4:0] inputBram_io_b_addr;
  wire [15:0] inputBram_io_b_dout;
  reg [4:0] inputReadAddr;
  reg [31:0] _RAND_37;
  reg  inputPieceRead;
  reg [31:0] _RAND_38;
  wire  outputBram_clock;
  wire [4:0] outputBram_io_a_addr;
  wire [15:0] outputBram_io_a_din;
  wire  outputBram_io_a_wr;
  wire [4:0] outputBram_io_b_addr;
  wire [15:0] outputBram_io_b_dout;
  reg [4:0] outputWriteAddr;
  reg [31:0] _RAND_39;
  reg [4:0] outputReadAddr;
  reg [31:0] _RAND_40;
  wire  _T_75;
  wire  _T_76;
  wire  _GEN_0;
  wire [9:0] _GEN_1;
  wire  _T_79;
  wire  _T_80;
  wire  _GEN_2;
  wire  _T_84;
  wire  _T_85;
  wire  _T_87;
  wire  _T_88;
  wire  _T_90;
  wire  _T_94;
  wire [9:0] _T_96;
  wire [5:0] _T_98;
  wire [4:0] _T_99;
  wire  _T_100;
  wire  _T_101;
  wire  _T_102;
  wire  _T_103;
  wire  _T_104;
  wire  _T_105;
  wire  _T_106;
  wire  _T_107;
  wire  _T_108;
  wire  _T_109;
  wire  _T_110;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  _T_114;
  wire  _T_115;
  wire [9:0] _GEN_4;
  wire [4:0] _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [9:0] _GEN_23;
  wire [4:0] _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  inputAdvance;
  wire  _T_118;
  wire  _T_120;
  wire  _T_122;
  wire  _T_123;
  wire  _T_125;
  wire  _T_126;
  wire [5:0] _T_128;
  wire [5:0] _T_129;
  wire [4:0] _T_130;
  wire [10:0] _T_132;
  wire [10:0] _T_133;
  wire [9:0] _T_134;
  wire [9:0] _GEN_41;
  wire [9:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  nextBitValid;
  wire  nextBit;
  wire [5:0] _T_138;
  wire [4:0] _T_139;
  wire [10:0] _T_141;
  wire [9:0] _T_142;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire [4:0] _GEN_74;
  wire [9:0] _GEN_75;
  wire  _T_144;
  wire  _T_147;
  wire  _T_149;
  wire  _T_150;
  wire  _T_151;
  wire [1:0] _T_152;
  wire [1:0] _T_153;
  wire [3:0] _T_154;
  wire [1:0] _T_155;
  wire [1:0] _T_156;
  wire [3:0] _T_157;
  wire [7:0] _T_158;
  wire [1:0] _T_159;
  wire [1:0] _T_160;
  wire [3:0] _T_161;
  wire [1:0] _T_162;
  wire [1:0] _T_163;
  wire [3:0] _T_164;
  wire [7:0] _T_165;
  wire [15:0] _T_166;
  wire [5:0] _T_171;
  wire [4:0] _T_172;
  wire [4:0] _GEN_76;
  wire [4:0] _GEN_77;
  reg  outputReadingStarted;
  reg [31:0] _RAND_41;
  wire  _T_177;
  wire  _T_184;
  wire  _T_185;
  wire  _T_186;
  wire  _T_187;
  wire  _GEN_78;
  wire  _T_189;
  wire  _T_191;
  wire  _T_192;
  wire [5:0] _T_194;
  wire [4:0] _T_195;
  wire [4:0] _GEN_79;
  wire  _T_199;
  wire  _T_200;
  wire  _T_210;
  wire  _T_215;
  wire  _T_216;
  wire [9:0] _GEN_80;
  wire [4:0] _GEN_81;
  wire  _GEN_82;
  wire [4:0] _GEN_83;
  wire [4:0] _GEN_84;
  DualPortBRAM inputBram (
    .clock(inputBram_clock),
    .io_a_addr(inputBram_io_a_addr),
    .io_a_din(inputBram_io_a_din),
    .io_a_wr(inputBram_io_a_wr),
    .io_b_addr(inputBram_io_b_addr),
    .io_b_dout(inputBram_io_b_dout)
  );
  DualPortBRAM outputBram (
    .clock(outputBram_clock),
    .io_a_addr(outputBram_io_a_addr),
    .io_a_din(outputBram_io_a_din),
    .io_a_wr(outputBram_io_a_wr),
    .io_b_addr(outputBram_io_b_addr),
    .io_b_dout(outputBram_io_b_dout)
  );
  assign _T_75 = io_inputMemIdx == 5'h1f;
  assign _T_76 = io_inputMemBlockValid & _T_75;
  assign _GEN_0 = _T_76 ? 1'h1 : inputBlockLoaded;
  assign _GEN_1 = _T_76 ? io_inputBits : inputBitsRemaining;
  assign _T_79 = inputBitsRemaining == 10'h0;
  assign _T_80 = inputBlockLoaded & _T_79;
  assign _GEN_2 = _T_80 ? 1'h0 : _GEN_0;
  assign _T_84 = inputPieceBitsRemaining == 5'h0;
  assign _T_85 = inputBlockLoaded & _T_84;
  assign _T_87 = inputBitsRemaining != 10'h0;
  assign _T_88 = _T_85 & _T_87;
  assign _T_90 = inputPieceRead == 1'h0;
  assign _T_94 = inputBitsRemaining < 10'h10;
  assign _T_96 = _T_94 ? inputBitsRemaining : 10'h10;
  assign _T_98 = inputReadAddr + 5'h1;
  assign _T_99 = _T_98[4:0];
  assign _T_100 = inputBram_io_b_dout[0];
  assign _T_101 = inputBram_io_b_dout[1];
  assign _T_102 = inputBram_io_b_dout[2];
  assign _T_103 = inputBram_io_b_dout[3];
  assign _T_104 = inputBram_io_b_dout[4];
  assign _T_105 = inputBram_io_b_dout[5];
  assign _T_106 = inputBram_io_b_dout[6];
  assign _T_107 = inputBram_io_b_dout[7];
  assign _T_108 = inputBram_io_b_dout[8];
  assign _T_109 = inputBram_io_b_dout[9];
  assign _T_110 = inputBram_io_b_dout[10];
  assign _T_111 = inputBram_io_b_dout[11];
  assign _T_112 = inputBram_io_b_dout[12];
  assign _T_113 = inputBram_io_b_dout[13];
  assign _T_114 = inputBram_io_b_dout[14];
  assign _T_115 = inputBram_io_b_dout[15];
  assign _GEN_4 = _T_90 ? {{5'd0}, inputPieceBitsRemaining} : _T_96;
  assign _GEN_5 = _T_90 ? inputReadAddr : _T_99;
  assign _GEN_6 = _T_90 ? inputMemBlock_0 : _T_100;
  assign _GEN_7 = _T_90 ? inputMemBlock_1 : _T_101;
  assign _GEN_8 = _T_90 ? inputMemBlock_2 : _T_102;
  assign _GEN_9 = _T_90 ? inputMemBlock_3 : _T_103;
  assign _GEN_10 = _T_90 ? inputMemBlock_4 : _T_104;
  assign _GEN_11 = _T_90 ? inputMemBlock_5 : _T_105;
  assign _GEN_12 = _T_90 ? inputMemBlock_6 : _T_106;
  assign _GEN_13 = _T_90 ? inputMemBlock_7 : _T_107;
  assign _GEN_14 = _T_90 ? inputMemBlock_8 : _T_108;
  assign _GEN_15 = _T_90 ? inputMemBlock_9 : _T_109;
  assign _GEN_16 = _T_90 ? inputMemBlock_10 : _T_110;
  assign _GEN_17 = _T_90 ? inputMemBlock_11 : _T_111;
  assign _GEN_18 = _T_90 ? inputMemBlock_12 : _T_112;
  assign _GEN_19 = _T_90 ? inputMemBlock_13 : _T_113;
  assign _GEN_20 = _T_90 ? inputMemBlock_14 : _T_114;
  assign _GEN_21 = _T_90 ? inputMemBlock_15 : _T_115;
  assign _GEN_22 = _T_88 ? _T_90 : inputPieceRead;
  assign _GEN_23 = _T_88 ? _GEN_4 : {{5'd0}, inputPieceBitsRemaining};
  assign _GEN_24 = _T_88 ? _GEN_5 : inputReadAddr;
  assign _GEN_25 = _T_88 ? _GEN_6 : inputMemBlock_0;
  assign _GEN_26 = _T_88 ? _GEN_7 : inputMemBlock_1;
  assign _GEN_27 = _T_88 ? _GEN_8 : inputMemBlock_2;
  assign _GEN_28 = _T_88 ? _GEN_9 : inputMemBlock_3;
  assign _GEN_29 = _T_88 ? _GEN_10 : inputMemBlock_4;
  assign _GEN_30 = _T_88 ? _GEN_11 : inputMemBlock_5;
  assign _GEN_31 = _T_88 ? _GEN_12 : inputMemBlock_6;
  assign _GEN_32 = _T_88 ? _GEN_13 : inputMemBlock_7;
  assign _GEN_33 = _T_88 ? _GEN_14 : inputMemBlock_8;
  assign _GEN_34 = _T_88 ? _GEN_15 : inputMemBlock_9;
  assign _GEN_35 = _T_88 ? _GEN_16 : inputMemBlock_10;
  assign _GEN_36 = _T_88 ? _GEN_17 : inputMemBlock_11;
  assign _GEN_37 = _T_88 ? _GEN_18 : inputMemBlock_12;
  assign _GEN_38 = _T_88 ? _GEN_19 : inputMemBlock_13;
  assign _GEN_39 = _T_88 ? _GEN_20 : inputMemBlock_14;
  assign _GEN_40 = _T_88 ? _GEN_21 : inputMemBlock_15;
  assign _T_118 = outputPieceBits != 5'h10;
  assign _T_120 = outputBits == 10'h200;
  assign _T_122 = _T_120 == 1'h0;
  assign _T_123 = _T_118 & _T_122;
  assign _T_125 = inputPieceBitsRemaining != 5'h0;
  assign _T_126 = _T_123 & _T_125;
  assign _T_128 = inputPieceBitsRemaining - 5'h1;
  assign _T_129 = $unsigned(_T_128);
  assign _T_130 = _T_129[4:0];
  assign _T_132 = inputBitsRemaining - 10'h1;
  assign _T_133 = $unsigned(_T_132);
  assign _T_134 = _T_133[9:0];
  assign _GEN_41 = inputAdvance ? {{5'd0}, _T_130} : _GEN_23;
  assign _GEN_42 = inputAdvance ? _T_134 : _GEN_1;
  assign _GEN_43 = inputAdvance ? inputMemBlock_1 : _GEN_25;
  assign _GEN_44 = inputAdvance ? inputMemBlock_2 : _GEN_26;
  assign _GEN_45 = inputAdvance ? inputMemBlock_3 : _GEN_27;
  assign _GEN_46 = inputAdvance ? inputMemBlock_4 : _GEN_28;
  assign _GEN_47 = inputAdvance ? inputMemBlock_5 : _GEN_29;
  assign _GEN_48 = inputAdvance ? inputMemBlock_6 : _GEN_30;
  assign _GEN_49 = inputAdvance ? inputMemBlock_7 : _GEN_31;
  assign _GEN_50 = inputAdvance ? inputMemBlock_8 : _GEN_32;
  assign _GEN_51 = inputAdvance ? inputMemBlock_9 : _GEN_33;
  assign _GEN_52 = inputAdvance ? inputMemBlock_10 : _GEN_34;
  assign _GEN_53 = inputAdvance ? inputMemBlock_11 : _GEN_35;
  assign _GEN_54 = inputAdvance ? inputMemBlock_12 : _GEN_36;
  assign _GEN_55 = inputAdvance ? inputMemBlock_13 : _GEN_37;
  assign _GEN_56 = inputAdvance ? inputMemBlock_14 : _GEN_38;
  assign _GEN_57 = inputAdvance ? inputMemBlock_15 : _GEN_39;
  assign _T_138 = outputPieceBits + 5'h1;
  assign _T_139 = _T_138[4:0];
  assign _T_141 = outputBits + 10'h1;
  assign _T_142 = _T_141[9:0];
  assign _GEN_58 = nextBitValid ? nextBit : outputMemBlock_15;
  assign _GEN_59 = nextBitValid ? outputMemBlock_1 : outputMemBlock_0;
  assign _GEN_60 = nextBitValid ? outputMemBlock_2 : outputMemBlock_1;
  assign _GEN_61 = nextBitValid ? outputMemBlock_3 : outputMemBlock_2;
  assign _GEN_62 = nextBitValid ? outputMemBlock_4 : outputMemBlock_3;
  assign _GEN_63 = nextBitValid ? outputMemBlock_5 : outputMemBlock_4;
  assign _GEN_64 = nextBitValid ? outputMemBlock_6 : outputMemBlock_5;
  assign _GEN_65 = nextBitValid ? outputMemBlock_7 : outputMemBlock_6;
  assign _GEN_66 = nextBitValid ? outputMemBlock_8 : outputMemBlock_7;
  assign _GEN_67 = nextBitValid ? outputMemBlock_9 : outputMemBlock_8;
  assign _GEN_68 = nextBitValid ? outputMemBlock_10 : outputMemBlock_9;
  assign _GEN_69 = nextBitValid ? outputMemBlock_11 : outputMemBlock_10;
  assign _GEN_70 = nextBitValid ? outputMemBlock_12 : outputMemBlock_11;
  assign _GEN_71 = nextBitValid ? outputMemBlock_13 : outputMemBlock_12;
  assign _GEN_72 = nextBitValid ? outputMemBlock_14 : outputMemBlock_13;
  assign _GEN_73 = nextBitValid ? outputMemBlock_15 : outputMemBlock_14;
  assign _GEN_74 = nextBitValid ? _T_139 : outputPieceBits;
  assign _GEN_75 = nextBitValid ? _T_142 : outputBits;
  assign _T_144 = outputPieceBits == 5'h10;
  assign _T_147 = io_inputFinished & _T_79;
  assign _T_149 = outputPieceBits > 5'h0;
  assign _T_150 = _T_147 & _T_149;
  assign _T_151 = _T_144 | _T_150;
  assign _T_152 = {outputMemBlock_1,outputMemBlock_0};
  assign _T_153 = {outputMemBlock_3,outputMemBlock_2};
  assign _T_154 = {_T_153,_T_152};
  assign _T_155 = {outputMemBlock_5,outputMemBlock_4};
  assign _T_156 = {outputMemBlock_7,outputMemBlock_6};
  assign _T_157 = {_T_156,_T_155};
  assign _T_158 = {_T_157,_T_154};
  assign _T_159 = {outputMemBlock_9,outputMemBlock_8};
  assign _T_160 = {outputMemBlock_11,outputMemBlock_10};
  assign _T_161 = {_T_160,_T_159};
  assign _T_162 = {outputMemBlock_13,outputMemBlock_12};
  assign _T_163 = {outputMemBlock_15,outputMemBlock_14};
  assign _T_164 = {_T_163,_T_162};
  assign _T_165 = {_T_164,_T_161};
  assign _T_166 = {_T_165,_T_158};
  assign _T_171 = outputWriteAddr + 5'h1;
  assign _T_172 = _T_171[4:0];
  assign _GEN_76 = _T_144 ? 5'h0 : _GEN_74;
  assign _GEN_77 = _T_144 ? _T_172 : outputWriteAddr;
  assign _T_177 = outputReadingStarted == 1'h0;
  assign _T_184 = outputBits > 10'h0;
  assign _T_185 = _T_147 & _T_184;
  assign _T_186 = _T_120 | _T_185;
  assign _T_187 = _T_177 & _T_186;
  assign _GEN_78 = _T_187 ? 1'h1 : outputReadingStarted;
  assign _T_189 = io_outputMemBlockReady & outputReadingStarted;
  assign _T_191 = outputReadAddr != 5'h1f;
  assign _T_192 = _T_189 & _T_191;
  assign _T_194 = outputReadAddr + 5'h1;
  assign _T_195 = _T_194[4:0];
  assign _GEN_79 = _T_192 ? _T_195 : outputReadAddr;
  assign _T_199 = io_inputFinished == 1'h0;
  assign _T_200 = _T_79 & _T_199;
  assign _T_210 = outputReadingStarted & _T_186;
  assign _T_215 = outputBits == 10'h0;
  assign _T_216 = _T_147 & _T_215;
  assign _GEN_80 = io_outputMemFlushed ? 10'h0 : _GEN_75;
  assign _GEN_81 = io_outputMemFlushed ? 5'h0 : _GEN_76;
  assign _GEN_82 = io_outputMemFlushed ? 1'h0 : _GEN_78;
  assign _GEN_83 = io_outputMemFlushed ? 5'h0 : _GEN_77;
  assign _GEN_84 = io_outputMemFlushed ? 5'h0 : _GEN_79;
  assign io_inputMemConsumed = _T_200;
  assign io_outputMemBlock = outputBram_io_b_dout;
  assign io_outputMemBlockValid = _T_210;
  assign io_outputBits = outputBits;
  assign io_outputFinished = _T_216;
  assign inputBram_io_a_addr = io_inputMemIdx;
  assign inputBram_io_a_din = io_inputMemBlock;
  assign inputBram_io_a_wr = io_inputMemBlockValid;
  assign inputBram_io_b_addr = inputReadAddr;
  assign inputBram_clock = clock;
  assign outputBram_io_a_addr = outputWriteAddr;
  assign outputBram_io_a_din = _T_166;
  assign outputBram_io_a_wr = _T_151;
  assign outputBram_io_b_addr = outputReadAddr;
  assign outputBram_clock = clock;
  assign inputAdvance = _T_126;
  assign nextBitValid = inputAdvance;
  assign nextBit = inputMemBlock_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  inputMemBlock_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  inputMemBlock_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputMemBlock_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  inputMemBlock_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  inputMemBlock_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  inputMemBlock_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  inputMemBlock_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemBlock_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBlock_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  inputMemBlock_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputMemBlock_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  inputMemBlock_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  inputMemBlock_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  inputMemBlock_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  inputMemBlock_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  inputMemBlock_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  inputPieceBitsRemaining = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  inputBitsRemaining = _RAND_17[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  inputBlockLoaded = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  outputMemBlock_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  outputMemBlock_1 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  outputMemBlock_2 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  outputMemBlock_3 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  outputMemBlock_4 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  outputMemBlock_5 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  outputMemBlock_6 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  outputMemBlock_7 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  outputMemBlock_8 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  outputMemBlock_9 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  outputMemBlock_10 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  outputMemBlock_11 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  outputMemBlock_12 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  outputMemBlock_13 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  outputMemBlock_14 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  outputMemBlock_15 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  outputBits = _RAND_35[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  outputPieceBits = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  inputReadAddr = _RAND_37[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  inputPieceRead = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  outputWriteAddr = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  outputReadAddr = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  outputReadingStarted = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (inputAdvance) begin
      inputMemBlock_0 <= inputMemBlock_1;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_0 <= _T_100;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_1 <= inputMemBlock_2;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_1 <= _T_101;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_2 <= inputMemBlock_3;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_2 <= _T_102;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_3 <= inputMemBlock_4;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_3 <= _T_103;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_4 <= inputMemBlock_5;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_4 <= _T_104;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_5 <= inputMemBlock_6;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_5 <= _T_105;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_6 <= inputMemBlock_7;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_6 <= _T_106;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_7 <= inputMemBlock_8;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_7 <= _T_107;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_8 <= inputMemBlock_9;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_8 <= _T_108;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_9 <= inputMemBlock_10;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_9 <= _T_109;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_10 <= inputMemBlock_11;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_10 <= _T_110;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_11 <= inputMemBlock_12;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_11 <= _T_111;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_12 <= inputMemBlock_13;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_12 <= _T_112;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_13 <= inputMemBlock_14;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_13 <= _T_113;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_14 <= inputMemBlock_15;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputMemBlock_14 <= _T_114;
        end
      end
    end
    if (_T_88) begin
      if (!(_T_90)) begin
        inputMemBlock_15 <= _T_115;
      end
    end
    if (reset) begin
      inputPieceBitsRemaining <= 5'h0;
    end else begin
      inputPieceBitsRemaining <= _GEN_41[4:0];
    end
    if (reset) begin
      inputBitsRemaining <= 10'h0;
    end else begin
      if (inputAdvance) begin
        inputBitsRemaining <= _T_134;
      end else begin
        if (_T_76) begin
          inputBitsRemaining <= io_inputBits;
        end
      end
    end
    if (reset) begin
      inputBlockLoaded <= 1'h0;
    end else begin
      if (_T_80) begin
        inputBlockLoaded <= 1'h0;
      end else begin
        if (_T_76) begin
          inputBlockLoaded <= 1'h1;
        end
      end
    end
    if (nextBitValid) begin
      outputMemBlock_0 <= outputMemBlock_1;
    end
    if (nextBitValid) begin
      outputMemBlock_1 <= outputMemBlock_2;
    end
    if (nextBitValid) begin
      outputMemBlock_2 <= outputMemBlock_3;
    end
    if (nextBitValid) begin
      outputMemBlock_3 <= outputMemBlock_4;
    end
    if (nextBitValid) begin
      outputMemBlock_4 <= outputMemBlock_5;
    end
    if (nextBitValid) begin
      outputMemBlock_5 <= outputMemBlock_6;
    end
    if (nextBitValid) begin
      outputMemBlock_6 <= outputMemBlock_7;
    end
    if (nextBitValid) begin
      outputMemBlock_7 <= outputMemBlock_8;
    end
    if (nextBitValid) begin
      outputMemBlock_8 <= outputMemBlock_9;
    end
    if (nextBitValid) begin
      outputMemBlock_9 <= outputMemBlock_10;
    end
    if (nextBitValid) begin
      outputMemBlock_10 <= outputMemBlock_11;
    end
    if (nextBitValid) begin
      outputMemBlock_11 <= outputMemBlock_12;
    end
    if (nextBitValid) begin
      outputMemBlock_12 <= outputMemBlock_13;
    end
    if (nextBitValid) begin
      outputMemBlock_13 <= outputMemBlock_14;
    end
    if (nextBitValid) begin
      outputMemBlock_14 <= outputMemBlock_15;
    end
    if (nextBitValid) begin
      outputMemBlock_15 <= nextBit;
    end
    if (reset) begin
      outputBits <= 10'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputBits <= 10'h0;
      end else begin
        if (nextBitValid) begin
          outputBits <= _T_142;
        end
      end
    end
    if (reset) begin
      outputPieceBits <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputPieceBits <= 5'h0;
      end else begin
        if (_T_144) begin
          outputPieceBits <= 5'h0;
        end else begin
          if (nextBitValid) begin
            outputPieceBits <= _T_139;
          end
        end
      end
    end
    if (reset) begin
      inputReadAddr <= 5'h0;
    end else begin
      if (_T_88) begin
        if (!(_T_90)) begin
          inputReadAddr <= _T_99;
        end
      end
    end
    if (reset) begin
      inputPieceRead <= 1'h0;
    end else begin
      if (_T_88) begin
        inputPieceRead <= _T_90;
      end
    end
    if (reset) begin
      outputWriteAddr <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputWriteAddr <= 5'h0;
      end else begin
        if (_T_144) begin
          outputWriteAddr <= _T_172;
        end
      end
    end
    if (reset) begin
      outputReadAddr <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputReadAddr <= 5'h0;
      end else begin
        if (_T_192) begin
          outputReadAddr <= _T_195;
        end
      end
    end
    if (reset) begin
      outputReadingStarted <= 1'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputReadingStarted <= 1'h0;
      end else begin
        if (_T_187) begin
          outputReadingStarted <= 1'h1;
        end
      end
    end
  end
endmodule
module StreamingCore(
  input         clock,
  input         reset,
  output [63:0] io_inputMemAddr,
  output        io_inputMemAddrValid,
  input         io_inputMemAddrReady,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output        io_inputMemBlockReady,
  output [63:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [15:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output        io_inputFinished,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [15:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [15:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [63:0] inputBitsRemaining;
  reg [63:0] _RAND_2;
  reg  coreInputFinished;
  reg [31:0] _RAND_3;
  reg [63:0] outputBits;
  reg [63:0] _RAND_4;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_5;
  reg  outputLengthCommitted;
  reg [31:0] _RAND_6;
  reg [63:0] inputMemAddr;
  reg [63:0] _RAND_7;
  reg [63:0] outputMemAddr;
  reg [63:0] _RAND_8;
  reg [63:0] outputLenAddr;
  reg [63:0] _RAND_9;
  reg  inputAddressAccepted;
  reg [31:0] _RAND_10;
  wire  _T_41;
  wire  _T_42;
  wire  _T_44;
  wire  _T_46;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_53;
  wire  _GEN_0;
  wire  inputBlockReadable;
  wire  _T_56;
  wire  _T_57;
  wire  _T_59;
  wire [9:0] _T_61;
  wire [9:0] _T_62;
  wire  _T_64;
  wire [47:0] _T_65;
  wire [63:0] _T_66;
  wire [63:0] _GEN_1;
  wire  _T_68;
  wire [31:0] _T_69;
  wire [47:0] _T_70;
  wire [15:0] _T_71;
  wire [63:0] _T_72;
  wire [63:0] _GEN_2;
  wire  _T_74;
  wire [15:0] _T_75;
  wire [31:0] _T_76;
  wire [31:0] _T_77;
  wire [63:0] _T_78;
  wire [63:0] _GEN_3;
  wire  _T_80;
  wire [47:0] _T_81;
  wire [63:0] _T_82;
  wire [63:0] _GEN_4;
  wire  _T_84;
  wire [47:0] _T_85;
  wire [63:0] _T_86;
  wire [63:0] _GEN_5;
  wire  _T_88;
  wire [31:0] _T_89;
  wire [47:0] _T_90;
  wire [15:0] _T_91;
  wire [63:0] _T_92;
  wire [63:0] _GEN_6;
  wire  _T_94;
  wire [15:0] _T_95;
  wire [31:0] _T_96;
  wire [31:0] _T_97;
  wire [63:0] _T_98;
  wire [63:0] _GEN_7;
  wire  _T_100;
  wire [47:0] _T_101;
  wire [63:0] _T_102;
  wire [63:0] _GEN_8;
  wire  _T_104;
  wire [47:0] _T_105;
  wire [63:0] _T_106;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire  _T_108;
  wire [31:0] _T_109;
  wire [47:0] _T_110;
  wire [15:0] _T_111;
  wire [63:0] _T_112;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire  _T_114;
  wire [15:0] _T_115;
  wire [31:0] _T_116;
  wire [31:0] _T_117;
  wire [63:0] _T_118;
  wire [63:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire  _T_120;
  wire [47:0] _T_121;
  wire [63:0] _T_122;
  wire [63:0] _GEN_15;
  wire [63:0] _GEN_16;
  wire  _T_124;
  wire [64:0] _T_128;
  wire [63:0] _T_129;
  wire  _GEN_17;
  wire  _GEN_18;
  wire [63:0] _GEN_19;
  wire [64:0] _T_135;
  wire [64:0] _T_136;
  wire [63:0] _T_137;
  wire [63:0] _T_139;
  wire [64:0] _T_141;
  wire [63:0] _T_142;
  wire [63:0] _GEN_20;
  wire [63:0] _GEN_21;
  wire [63:0] _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [63:0] _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire [63:0] _GEN_29;
  wire [63:0] _GEN_30;
  wire [63:0] _GEN_31;
  wire [63:0] _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _T_150;
  wire  _GEN_36;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_11;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_12;
  wire  _GEN_37;
  wire [63:0] _T_157;
  wire  _T_159;
  wire  _T_161;
  wire  _T_162;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _GEN_38;
  wire  _T_171;
  wire [4:0] _GEN_39;
  wire [5:0] _T_174;
  wire [4:0] _T_175;
  wire [4:0] _GEN_40;
  wire [4:0] _GEN_41;
  wire [15:0] outputBitsBlock;
  wire  _T_178;
  wire [15:0] _T_179;
  wire  _T_181;
  wire [15:0] _T_182;
  wire  _T_184;
  wire [15:0] _T_185;
  wire  _T_187;
  wire [15:0] _T_188;
  wire [15:0] _T_190;
  wire [15:0] _T_191;
  wire [15:0] _T_192;
  wire [15:0] _T_193;
  wire [15:0] _T_194;
  wire  _T_195;
  wire  _T_199;
  wire [63:0] _GEN_50;
  wire [64:0] _T_203;
  wire [63:0] _T_204;
  wire  _GEN_42;
  wire [63:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire [63:0] _GEN_48;
  wire [63:0] _GEN_49;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign _T_41 = inputAddressAccepted == 1'h0;
  assign _T_42 = initDone & core_io_inputMemConsumed;
  assign _T_44 = inputBitsRemaining == 64'h0;
  assign _T_46 = _T_44 == 1'h0;
  assign _T_47 = _T_42 & _T_46;
  assign _T_48 = isInit | _T_47;
  assign _T_49 = _T_41 & _T_48;
  assign _T_50 = io_inputMemAddrValid & io_inputMemAddrReady;
  assign _T_53 = reset == 1'h0;
  assign _GEN_0 = _T_50 ? 1'h1 : inputAddressAccepted;
  assign _T_56 = inputAddressAccepted & io_inputMemBlockValid;
  assign _T_57 = inputBlockReadable & initDone;
  assign _T_59 = inputBitsRemaining > 64'h200;
  assign _T_61 = inputBitsRemaining[9:0];
  assign _T_62 = _T_59 ? 10'h200 : _T_61;
  assign _T_64 = io_inputMemIdx == 5'h0;
  assign _T_65 = inputMemAddr[63:16];
  assign _T_66 = {_T_65,io_inputMemBlock};
  assign _GEN_1 = _T_64 ? _T_66 : inputMemAddr;
  assign _T_68 = io_inputMemIdx == 5'h1;
  assign _T_69 = inputMemAddr[63:32];
  assign _T_70 = {_T_69,io_inputMemBlock};
  assign _T_71 = inputMemAddr[15:0];
  assign _T_72 = {_T_70,_T_71};
  assign _GEN_2 = _T_68 ? _T_72 : _GEN_1;
  assign _T_74 = io_inputMemIdx == 5'h2;
  assign _T_75 = inputMemAddr[63:48];
  assign _T_76 = {_T_75,io_inputMemBlock};
  assign _T_77 = inputMemAddr[31:0];
  assign _T_78 = {_T_76,_T_77};
  assign _GEN_3 = _T_74 ? _T_78 : _GEN_2;
  assign _T_80 = io_inputMemIdx == 5'h3;
  assign _T_81 = inputMemAddr[47:0];
  assign _T_82 = {io_inputMemBlock,_T_81};
  assign _GEN_4 = _T_80 ? _T_82 : _GEN_3;
  assign _T_84 = io_inputMemIdx == 5'h4;
  assign _T_85 = inputBitsRemaining[63:16];
  assign _T_86 = {_T_85,io_inputMemBlock};
  assign _GEN_5 = _T_84 ? _T_86 : inputBitsRemaining;
  assign _T_88 = io_inputMemIdx == 5'h5;
  assign _T_89 = inputBitsRemaining[63:32];
  assign _T_90 = {_T_89,io_inputMemBlock};
  assign _T_91 = inputBitsRemaining[15:0];
  assign _T_92 = {_T_90,_T_91};
  assign _GEN_6 = _T_88 ? _T_92 : _GEN_5;
  assign _T_94 = io_inputMemIdx == 5'h6;
  assign _T_95 = inputBitsRemaining[63:48];
  assign _T_96 = {_T_95,io_inputMemBlock};
  assign _T_97 = inputBitsRemaining[31:0];
  assign _T_98 = {_T_96,_T_97};
  assign _GEN_7 = _T_94 ? _T_98 : _GEN_6;
  assign _T_100 = io_inputMemIdx == 5'h7;
  assign _T_101 = inputBitsRemaining[47:0];
  assign _T_102 = {io_inputMemBlock,_T_101};
  assign _GEN_8 = _T_100 ? _T_102 : _GEN_7;
  assign _T_104 = io_inputMemIdx == 5'h8;
  assign _T_105 = outputMemAddr[63:16];
  assign _T_106 = {_T_105,io_inputMemBlock};
  assign _GEN_9 = _T_104 ? _T_106 : outputMemAddr;
  assign _GEN_10 = _T_104 ? _T_106 : outputLenAddr;
  assign _T_108 = io_inputMemIdx == 5'h9;
  assign _T_109 = outputMemAddr[63:32];
  assign _T_110 = {_T_109,io_inputMemBlock};
  assign _T_111 = outputMemAddr[15:0];
  assign _T_112 = {_T_110,_T_111};
  assign _GEN_11 = _T_108 ? _T_112 : _GEN_9;
  assign _GEN_12 = _T_108 ? _T_112 : _GEN_10;
  assign _T_114 = io_inputMemIdx == 5'ha;
  assign _T_115 = outputMemAddr[63:48];
  assign _T_116 = {_T_115,io_inputMemBlock};
  assign _T_117 = outputMemAddr[31:0];
  assign _T_118 = {_T_116,_T_117};
  assign _GEN_13 = _T_114 ? _T_118 : _GEN_11;
  assign _GEN_14 = _T_114 ? _T_118 : _GEN_12;
  assign _T_120 = io_inputMemIdx == 5'hb;
  assign _T_121 = outputMemAddr[47:0];
  assign _T_122 = {io_inputMemBlock,_T_121};
  assign _GEN_15 = _T_120 ? _T_122 : _GEN_13;
  assign _GEN_16 = _T_120 ? _T_122 : _GEN_14;
  assign _T_124 = io_inputMemIdx == 5'h1f;
  assign _T_128 = outputMemAddr + 64'h40;
  assign _T_129 = _T_128[63:0];
  assign _GEN_17 = _T_124 ? 1'h0 : isInit;
  assign _GEN_18 = _T_124 ? 1'h1 : initDone;
  assign _GEN_19 = _T_124 ? _T_129 : _GEN_15;
  assign _T_135 = inputBitsRemaining - 64'h200;
  assign _T_136 = $unsigned(_T_135);
  assign _T_137 = _T_136[63:0];
  assign _T_139 = _T_59 ? _T_137 : 64'h0;
  assign _T_141 = inputMemAddr + 64'h40;
  assign _T_142 = _T_141[63:0];
  assign _GEN_20 = _T_124 ? _T_139 : inputBitsRemaining;
  assign _GEN_21 = _T_124 ? _T_142 : inputMemAddr;
  assign _GEN_22 = isInit ? _GEN_4 : _GEN_21;
  assign _GEN_23 = isInit ? _GEN_8 : _GEN_20;
  assign _GEN_24 = isInit ? _GEN_19 : outputMemAddr;
  assign _GEN_25 = isInit ? _GEN_16 : outputLenAddr;
  assign _GEN_26 = isInit ? _GEN_17 : isInit;
  assign _GEN_27 = isInit ? _GEN_18 : initDone;
  assign _GEN_28 = _T_124 ? 1'h0 : _GEN_0;
  assign _GEN_29 = inputBlockReadable ? _GEN_22 : inputMemAddr;
  assign _GEN_30 = inputBlockReadable ? _GEN_23 : inputBitsRemaining;
  assign _GEN_31 = inputBlockReadable ? _GEN_24 : outputMemAddr;
  assign _GEN_32 = inputBlockReadable ? _GEN_25 : outputLenAddr;
  assign _GEN_33 = inputBlockReadable ? _GEN_26 : isInit;
  assign _GEN_34 = inputBlockReadable ? _GEN_27 : initDone;
  assign _GEN_35 = inputBlockReadable ? _GEN_28 : _GEN_0;
  assign _T_150 = core_io_inputMemConsumed & _T_44;
  assign _GEN_36 = _T_150 ? 1'h1 : coreInputFinished;
  assign _GEN_37 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_157 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_159 = outputAddressAccepted == 1'h0;
  assign _T_161 = outputLengthCommitted == 1'h0;
  assign _T_162 = core_io_outputFinished & _T_161;
  assign _T_163 = core_io_outputMemBlockValid | _T_162;
  assign _T_164 = _T_159 & _T_163;
  assign _T_165 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_38 = _T_165 ? 1'h1 : outputAddressAccepted;
  assign _T_171 = outputBlockCounter == 5'h1f;
  assign _GEN_39 = io_outputMemBlockReady ? 5'h0 : outputBlockCounter;
  assign _T_174 = outputBlockCounter + 5'h1;
  assign _T_175 = _T_174[4:0];
  assign _GEN_40 = _T_171 ? _GEN_39 : _T_175;
  assign _GEN_41 = outputAddressAcceptedNext ? _GEN_40 : outputBlockCounter;
  assign _T_178 = outputBlockCounter == 5'h0;
  assign _T_179 = outputBits[15:0];
  assign _T_181 = outputBlockCounter == 5'h1;
  assign _T_182 = outputBits[31:16];
  assign _T_184 = outputBlockCounter == 5'h2;
  assign _T_185 = outputBits[47:32];
  assign _T_187 = outputBlockCounter == 5'h3;
  assign _T_188 = outputBits[63:48];
  assign _T_190 = _T_187 ? _T_188 : 16'h0;
  assign _T_191 = _T_184 ? _T_185 : _T_190;
  assign _T_192 = _T_181 ? _T_182 : _T_191;
  assign _T_193 = _T_178 ? _T_179 : _T_192;
  assign _T_194 = core_io_outputFinished ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_195 = outputAddressAcceptedNext & io_outputMemBlockReady;
  assign _T_199 = _T_195 & _T_171;
  assign _GEN_50 = {{54'd0}, core_io_outputBits};
  assign _T_203 = outputBits + _GEN_50;
  assign _T_204 = _T_203[63:0];
  assign _GEN_42 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _GEN_43 = core_io_outputFinished ? outputBits : _T_204;
  assign _GEN_44 = core_io_outputFinished ? _GEN_31 : _T_129;
  assign _GEN_45 = _T_199 ? 1'h0 : _GEN_38;
  assign _GEN_46 = _T_199 ? 1'h0 : _GEN_37;
  assign _GEN_47 = _T_199 ? _GEN_42 : outputLengthCommitted;
  assign _GEN_48 = _T_199 ? _GEN_43 : outputBits;
  assign _GEN_49 = _T_199 ? _GEN_44 : _GEN_31;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemAddrValid = _T_49;
  assign io_inputMemBlockReady = inputAddressAccepted;
  assign io_outputMemAddr = _T_157;
  assign io_outputMemAddrValid = _T_164;
  assign io_outputMemBlock = _T_194;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_inputFinished = _T_44;
  assign io_outputFinished = outputLengthCommitted;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_57;
  assign core_io_inputBits = _T_62;
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_io_outputMemFlushed = _T_195;
  assign core_clock = clock;
  assign core_reset = reset;
  assign inputBlockReadable = _T_56;
  assign outputBitsBlock = _T_193;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{$random}};
  inputBitsRemaining = _RAND_2[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  coreInputFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{$random}};
  outputBits = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputBlockCounter = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputLengthCommitted = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{$random}};
  inputMemAddr = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{$random}};
  outputMemAddr = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{$random}};
  outputLenAddr = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputAddressAccepted = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  outputAddressAccepted = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  outputAddressAcceptedNext = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 64'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_100) begin
            inputBitsRemaining <= _T_102;
          end else begin
            if (_T_94) begin
              inputBitsRemaining <= _T_98;
            end else begin
              if (_T_88) begin
                inputBitsRemaining <= _T_92;
              end else begin
                if (_T_84) begin
                  inputBitsRemaining <= _T_86;
                end
              end
            end
          end
        end else begin
          if (_T_124) begin
            if (_T_59) begin
              inputBitsRemaining <= _T_137;
            end else begin
              inputBitsRemaining <= 64'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_150) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 64'h0;
    end else begin
      if (_T_199) begin
        if (!(core_io_outputFinished)) begin
          outputBits <= _T_204;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_171) begin
          if (io_outputMemBlockReady) begin
            outputBlockCounter <= 5'h0;
          end
        end else begin
          outputBlockCounter <= _T_175;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_199) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 64'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_80) begin
            inputMemAddr <= _T_82;
          end else begin
            if (_T_74) begin
              inputMemAddr <= _T_78;
            end else begin
              if (_T_68) begin
                inputMemAddr <= _T_72;
              end else begin
                if (_T_64) begin
                  inputMemAddr <= _T_66;
                end
              end
            end
          end
        end else begin
          if (_T_124) begin
            inputMemAddr <= _T_142;
          end
        end
      end
    end
    if (_T_199) begin
      if (core_io_outputFinished) begin
        if (inputBlockReadable) begin
          if (isInit) begin
            if (_T_124) begin
              outputMemAddr <= _T_129;
            end else begin
              if (_T_120) begin
                outputMemAddr <= _T_122;
              end else begin
                if (_T_114) begin
                  outputMemAddr <= _T_118;
                end else begin
                  if (_T_108) begin
                    outputMemAddr <= _T_112;
                  end else begin
                    if (_T_104) begin
                      outputMemAddr <= _T_106;
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        outputMemAddr <= _T_129;
      end
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            outputMemAddr <= _T_129;
          end else begin
            if (_T_120) begin
              outputMemAddr <= _T_122;
            end else begin
              if (_T_114) begin
                outputMemAddr <= _T_118;
              end else begin
                if (_T_108) begin
                  outputMemAddr <= _T_112;
                end else begin
                  if (_T_104) begin
                    outputMemAddr <= _T_106;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (inputBlockReadable) begin
      if (isInit) begin
        if (_T_120) begin
          outputLenAddr <= _T_122;
        end else begin
          if (_T_114) begin
            outputLenAddr <= _T_118;
          end else begin
            if (_T_108) begin
              outputLenAddr <= _T_112;
            end else begin
              if (_T_104) begin
                outputLenAddr <= _T_106;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      inputAddressAccepted <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (_T_124) begin
          inputAddressAccepted <= 1'h0;
        end else begin
          if (_T_50) begin
            inputAddressAccepted <= 1'h1;
          end
        end
      end else begin
        if (_T_50) begin
          inputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_199) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_165) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_199) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_50 & _T_53) begin
          $fwrite(32'h80000002,"input address 0x%h accepted for core 0\n",io_inputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_165 & _T_53) begin
          $fwrite(32'h80000002,"output address 0x%h accepted for core 0\n",io_outputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module StreamingCore_1(
  input         clock,
  input         reset,
  output [63:0] io_inputMemAddr,
  output        io_inputMemAddrValid,
  input         io_inputMemAddrReady,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output        io_inputMemBlockReady,
  output [63:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [15:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output        io_inputFinished,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [15:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [15:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [63:0] inputBitsRemaining;
  reg [63:0] _RAND_2;
  reg  coreInputFinished;
  reg [31:0] _RAND_3;
  reg [63:0] outputBits;
  reg [63:0] _RAND_4;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_5;
  reg  outputLengthCommitted;
  reg [31:0] _RAND_6;
  reg [63:0] inputMemAddr;
  reg [63:0] _RAND_7;
  reg [63:0] outputMemAddr;
  reg [63:0] _RAND_8;
  reg [63:0] outputLenAddr;
  reg [63:0] _RAND_9;
  reg  inputAddressAccepted;
  reg [31:0] _RAND_10;
  wire  _T_41;
  wire  _T_42;
  wire  _T_44;
  wire  _T_46;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_53;
  wire  _GEN_0;
  wire  inputBlockReadable;
  wire  _T_56;
  wire  _T_57;
  wire  _T_59;
  wire [9:0] _T_61;
  wire [9:0] _T_62;
  wire  _T_64;
  wire [47:0] _T_65;
  wire [63:0] _T_66;
  wire [63:0] _GEN_1;
  wire  _T_68;
  wire [31:0] _T_69;
  wire [47:0] _T_70;
  wire [15:0] _T_71;
  wire [63:0] _T_72;
  wire [63:0] _GEN_2;
  wire  _T_74;
  wire [15:0] _T_75;
  wire [31:0] _T_76;
  wire [31:0] _T_77;
  wire [63:0] _T_78;
  wire [63:0] _GEN_3;
  wire  _T_80;
  wire [47:0] _T_81;
  wire [63:0] _T_82;
  wire [63:0] _GEN_4;
  wire  _T_84;
  wire [47:0] _T_85;
  wire [63:0] _T_86;
  wire [63:0] _GEN_5;
  wire  _T_88;
  wire [31:0] _T_89;
  wire [47:0] _T_90;
  wire [15:0] _T_91;
  wire [63:0] _T_92;
  wire [63:0] _GEN_6;
  wire  _T_94;
  wire [15:0] _T_95;
  wire [31:0] _T_96;
  wire [31:0] _T_97;
  wire [63:0] _T_98;
  wire [63:0] _GEN_7;
  wire  _T_100;
  wire [47:0] _T_101;
  wire [63:0] _T_102;
  wire [63:0] _GEN_8;
  wire  _T_104;
  wire [47:0] _T_105;
  wire [63:0] _T_106;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire  _T_108;
  wire [31:0] _T_109;
  wire [47:0] _T_110;
  wire [15:0] _T_111;
  wire [63:0] _T_112;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire  _T_114;
  wire [15:0] _T_115;
  wire [31:0] _T_116;
  wire [31:0] _T_117;
  wire [63:0] _T_118;
  wire [63:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire  _T_120;
  wire [47:0] _T_121;
  wire [63:0] _T_122;
  wire [63:0] _GEN_15;
  wire [63:0] _GEN_16;
  wire  _T_124;
  wire [64:0] _T_128;
  wire [63:0] _T_129;
  wire  _GEN_17;
  wire  _GEN_18;
  wire [63:0] _GEN_19;
  wire [64:0] _T_135;
  wire [64:0] _T_136;
  wire [63:0] _T_137;
  wire [63:0] _T_139;
  wire [64:0] _T_141;
  wire [63:0] _T_142;
  wire [63:0] _GEN_20;
  wire [63:0] _GEN_21;
  wire [63:0] _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [63:0] _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire [63:0] _GEN_29;
  wire [63:0] _GEN_30;
  wire [63:0] _GEN_31;
  wire [63:0] _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _T_150;
  wire  _GEN_36;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_11;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_12;
  wire  _GEN_37;
  wire [63:0] _T_157;
  wire  _T_159;
  wire  _T_161;
  wire  _T_162;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _GEN_38;
  wire  _T_171;
  wire [4:0] _GEN_39;
  wire [5:0] _T_174;
  wire [4:0] _T_175;
  wire [4:0] _GEN_40;
  wire [4:0] _GEN_41;
  wire [15:0] outputBitsBlock;
  wire  _T_178;
  wire [15:0] _T_179;
  wire  _T_181;
  wire [15:0] _T_182;
  wire  _T_184;
  wire [15:0] _T_185;
  wire  _T_187;
  wire [15:0] _T_188;
  wire [15:0] _T_190;
  wire [15:0] _T_191;
  wire [15:0] _T_192;
  wire [15:0] _T_193;
  wire [15:0] _T_194;
  wire  _T_195;
  wire  _T_199;
  wire [63:0] _GEN_50;
  wire [64:0] _T_203;
  wire [63:0] _T_204;
  wire  _GEN_42;
  wire [63:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire [63:0] _GEN_48;
  wire [63:0] _GEN_49;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign _T_41 = inputAddressAccepted == 1'h0;
  assign _T_42 = initDone & core_io_inputMemConsumed;
  assign _T_44 = inputBitsRemaining == 64'h0;
  assign _T_46 = _T_44 == 1'h0;
  assign _T_47 = _T_42 & _T_46;
  assign _T_48 = isInit | _T_47;
  assign _T_49 = _T_41 & _T_48;
  assign _T_50 = io_inputMemAddrValid & io_inputMemAddrReady;
  assign _T_53 = reset == 1'h0;
  assign _GEN_0 = _T_50 ? 1'h1 : inputAddressAccepted;
  assign _T_56 = inputAddressAccepted & io_inputMemBlockValid;
  assign _T_57 = inputBlockReadable & initDone;
  assign _T_59 = inputBitsRemaining > 64'h200;
  assign _T_61 = inputBitsRemaining[9:0];
  assign _T_62 = _T_59 ? 10'h200 : _T_61;
  assign _T_64 = io_inputMemIdx == 5'h0;
  assign _T_65 = inputMemAddr[63:16];
  assign _T_66 = {_T_65,io_inputMemBlock};
  assign _GEN_1 = _T_64 ? _T_66 : inputMemAddr;
  assign _T_68 = io_inputMemIdx == 5'h1;
  assign _T_69 = inputMemAddr[63:32];
  assign _T_70 = {_T_69,io_inputMemBlock};
  assign _T_71 = inputMemAddr[15:0];
  assign _T_72 = {_T_70,_T_71};
  assign _GEN_2 = _T_68 ? _T_72 : _GEN_1;
  assign _T_74 = io_inputMemIdx == 5'h2;
  assign _T_75 = inputMemAddr[63:48];
  assign _T_76 = {_T_75,io_inputMemBlock};
  assign _T_77 = inputMemAddr[31:0];
  assign _T_78 = {_T_76,_T_77};
  assign _GEN_3 = _T_74 ? _T_78 : _GEN_2;
  assign _T_80 = io_inputMemIdx == 5'h3;
  assign _T_81 = inputMemAddr[47:0];
  assign _T_82 = {io_inputMemBlock,_T_81};
  assign _GEN_4 = _T_80 ? _T_82 : _GEN_3;
  assign _T_84 = io_inputMemIdx == 5'h4;
  assign _T_85 = inputBitsRemaining[63:16];
  assign _T_86 = {_T_85,io_inputMemBlock};
  assign _GEN_5 = _T_84 ? _T_86 : inputBitsRemaining;
  assign _T_88 = io_inputMemIdx == 5'h5;
  assign _T_89 = inputBitsRemaining[63:32];
  assign _T_90 = {_T_89,io_inputMemBlock};
  assign _T_91 = inputBitsRemaining[15:0];
  assign _T_92 = {_T_90,_T_91};
  assign _GEN_6 = _T_88 ? _T_92 : _GEN_5;
  assign _T_94 = io_inputMemIdx == 5'h6;
  assign _T_95 = inputBitsRemaining[63:48];
  assign _T_96 = {_T_95,io_inputMemBlock};
  assign _T_97 = inputBitsRemaining[31:0];
  assign _T_98 = {_T_96,_T_97};
  assign _GEN_7 = _T_94 ? _T_98 : _GEN_6;
  assign _T_100 = io_inputMemIdx == 5'h7;
  assign _T_101 = inputBitsRemaining[47:0];
  assign _T_102 = {io_inputMemBlock,_T_101};
  assign _GEN_8 = _T_100 ? _T_102 : _GEN_7;
  assign _T_104 = io_inputMemIdx == 5'h8;
  assign _T_105 = outputMemAddr[63:16];
  assign _T_106 = {_T_105,io_inputMemBlock};
  assign _GEN_9 = _T_104 ? _T_106 : outputMemAddr;
  assign _GEN_10 = _T_104 ? _T_106 : outputLenAddr;
  assign _T_108 = io_inputMemIdx == 5'h9;
  assign _T_109 = outputMemAddr[63:32];
  assign _T_110 = {_T_109,io_inputMemBlock};
  assign _T_111 = outputMemAddr[15:0];
  assign _T_112 = {_T_110,_T_111};
  assign _GEN_11 = _T_108 ? _T_112 : _GEN_9;
  assign _GEN_12 = _T_108 ? _T_112 : _GEN_10;
  assign _T_114 = io_inputMemIdx == 5'ha;
  assign _T_115 = outputMemAddr[63:48];
  assign _T_116 = {_T_115,io_inputMemBlock};
  assign _T_117 = outputMemAddr[31:0];
  assign _T_118 = {_T_116,_T_117};
  assign _GEN_13 = _T_114 ? _T_118 : _GEN_11;
  assign _GEN_14 = _T_114 ? _T_118 : _GEN_12;
  assign _T_120 = io_inputMemIdx == 5'hb;
  assign _T_121 = outputMemAddr[47:0];
  assign _T_122 = {io_inputMemBlock,_T_121};
  assign _GEN_15 = _T_120 ? _T_122 : _GEN_13;
  assign _GEN_16 = _T_120 ? _T_122 : _GEN_14;
  assign _T_124 = io_inputMemIdx == 5'h1f;
  assign _T_128 = outputMemAddr + 64'h40;
  assign _T_129 = _T_128[63:0];
  assign _GEN_17 = _T_124 ? 1'h0 : isInit;
  assign _GEN_18 = _T_124 ? 1'h1 : initDone;
  assign _GEN_19 = _T_124 ? _T_129 : _GEN_15;
  assign _T_135 = inputBitsRemaining - 64'h200;
  assign _T_136 = $unsigned(_T_135);
  assign _T_137 = _T_136[63:0];
  assign _T_139 = _T_59 ? _T_137 : 64'h0;
  assign _T_141 = inputMemAddr + 64'h40;
  assign _T_142 = _T_141[63:0];
  assign _GEN_20 = _T_124 ? _T_139 : inputBitsRemaining;
  assign _GEN_21 = _T_124 ? _T_142 : inputMemAddr;
  assign _GEN_22 = isInit ? _GEN_4 : _GEN_21;
  assign _GEN_23 = isInit ? _GEN_8 : _GEN_20;
  assign _GEN_24 = isInit ? _GEN_19 : outputMemAddr;
  assign _GEN_25 = isInit ? _GEN_16 : outputLenAddr;
  assign _GEN_26 = isInit ? _GEN_17 : isInit;
  assign _GEN_27 = isInit ? _GEN_18 : initDone;
  assign _GEN_28 = _T_124 ? 1'h0 : _GEN_0;
  assign _GEN_29 = inputBlockReadable ? _GEN_22 : inputMemAddr;
  assign _GEN_30 = inputBlockReadable ? _GEN_23 : inputBitsRemaining;
  assign _GEN_31 = inputBlockReadable ? _GEN_24 : outputMemAddr;
  assign _GEN_32 = inputBlockReadable ? _GEN_25 : outputLenAddr;
  assign _GEN_33 = inputBlockReadable ? _GEN_26 : isInit;
  assign _GEN_34 = inputBlockReadable ? _GEN_27 : initDone;
  assign _GEN_35 = inputBlockReadable ? _GEN_28 : _GEN_0;
  assign _T_150 = core_io_inputMemConsumed & _T_44;
  assign _GEN_36 = _T_150 ? 1'h1 : coreInputFinished;
  assign _GEN_37 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_157 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_159 = outputAddressAccepted == 1'h0;
  assign _T_161 = outputLengthCommitted == 1'h0;
  assign _T_162 = core_io_outputFinished & _T_161;
  assign _T_163 = core_io_outputMemBlockValid | _T_162;
  assign _T_164 = _T_159 & _T_163;
  assign _T_165 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_38 = _T_165 ? 1'h1 : outputAddressAccepted;
  assign _T_171 = outputBlockCounter == 5'h1f;
  assign _GEN_39 = io_outputMemBlockReady ? 5'h0 : outputBlockCounter;
  assign _T_174 = outputBlockCounter + 5'h1;
  assign _T_175 = _T_174[4:0];
  assign _GEN_40 = _T_171 ? _GEN_39 : _T_175;
  assign _GEN_41 = outputAddressAcceptedNext ? _GEN_40 : outputBlockCounter;
  assign _T_178 = outputBlockCounter == 5'h0;
  assign _T_179 = outputBits[15:0];
  assign _T_181 = outputBlockCounter == 5'h1;
  assign _T_182 = outputBits[31:16];
  assign _T_184 = outputBlockCounter == 5'h2;
  assign _T_185 = outputBits[47:32];
  assign _T_187 = outputBlockCounter == 5'h3;
  assign _T_188 = outputBits[63:48];
  assign _T_190 = _T_187 ? _T_188 : 16'h0;
  assign _T_191 = _T_184 ? _T_185 : _T_190;
  assign _T_192 = _T_181 ? _T_182 : _T_191;
  assign _T_193 = _T_178 ? _T_179 : _T_192;
  assign _T_194 = core_io_outputFinished ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_195 = outputAddressAcceptedNext & io_outputMemBlockReady;
  assign _T_199 = _T_195 & _T_171;
  assign _GEN_50 = {{54'd0}, core_io_outputBits};
  assign _T_203 = outputBits + _GEN_50;
  assign _T_204 = _T_203[63:0];
  assign _GEN_42 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _GEN_43 = core_io_outputFinished ? outputBits : _T_204;
  assign _GEN_44 = core_io_outputFinished ? _GEN_31 : _T_129;
  assign _GEN_45 = _T_199 ? 1'h0 : _GEN_38;
  assign _GEN_46 = _T_199 ? 1'h0 : _GEN_37;
  assign _GEN_47 = _T_199 ? _GEN_42 : outputLengthCommitted;
  assign _GEN_48 = _T_199 ? _GEN_43 : outputBits;
  assign _GEN_49 = _T_199 ? _GEN_44 : _GEN_31;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemAddrValid = _T_49;
  assign io_inputMemBlockReady = inputAddressAccepted;
  assign io_outputMemAddr = _T_157;
  assign io_outputMemAddrValid = _T_164;
  assign io_outputMemBlock = _T_194;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_inputFinished = _T_44;
  assign io_outputFinished = outputLengthCommitted;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_57;
  assign core_io_inputBits = _T_62;
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_io_outputMemFlushed = _T_195;
  assign core_clock = clock;
  assign core_reset = reset;
  assign inputBlockReadable = _T_56;
  assign outputBitsBlock = _T_193;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{$random}};
  inputBitsRemaining = _RAND_2[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  coreInputFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{$random}};
  outputBits = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputBlockCounter = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputLengthCommitted = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{$random}};
  inputMemAddr = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{$random}};
  outputMemAddr = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{$random}};
  outputLenAddr = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputAddressAccepted = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  outputAddressAccepted = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  outputAddressAcceptedNext = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 64'h1;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_100) begin
            inputBitsRemaining <= _T_102;
          end else begin
            if (_T_94) begin
              inputBitsRemaining <= _T_98;
            end else begin
              if (_T_88) begin
                inputBitsRemaining <= _T_92;
              end else begin
                if (_T_84) begin
                  inputBitsRemaining <= _T_86;
                end
              end
            end
          end
        end else begin
          if (_T_124) begin
            if (_T_59) begin
              inputBitsRemaining <= _T_137;
            end else begin
              inputBitsRemaining <= 64'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_150) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 64'h0;
    end else begin
      if (_T_199) begin
        if (!(core_io_outputFinished)) begin
          outputBits <= _T_204;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_171) begin
          if (io_outputMemBlockReady) begin
            outputBlockCounter <= 5'h0;
          end
        end else begin
          outputBlockCounter <= _T_175;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_199) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 64'h0;
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_80) begin
            inputMemAddr <= _T_82;
          end else begin
            if (_T_74) begin
              inputMemAddr <= _T_78;
            end else begin
              if (_T_68) begin
                inputMemAddr <= _T_72;
              end else begin
                if (_T_64) begin
                  inputMemAddr <= _T_66;
                end
              end
            end
          end
        end else begin
          if (_T_124) begin
            inputMemAddr <= _T_142;
          end
        end
      end
    end
    if (_T_199) begin
      if (core_io_outputFinished) begin
        if (inputBlockReadable) begin
          if (isInit) begin
            if (_T_124) begin
              outputMemAddr <= _T_129;
            end else begin
              if (_T_120) begin
                outputMemAddr <= _T_122;
              end else begin
                if (_T_114) begin
                  outputMemAddr <= _T_118;
                end else begin
                  if (_T_108) begin
                    outputMemAddr <= _T_112;
                  end else begin
                    if (_T_104) begin
                      outputMemAddr <= _T_106;
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        outputMemAddr <= _T_129;
      end
    end else begin
      if (inputBlockReadable) begin
        if (isInit) begin
          if (_T_124) begin
            outputMemAddr <= _T_129;
          end else begin
            if (_T_120) begin
              outputMemAddr <= _T_122;
            end else begin
              if (_T_114) begin
                outputMemAddr <= _T_118;
              end else begin
                if (_T_108) begin
                  outputMemAddr <= _T_112;
                end else begin
                  if (_T_104) begin
                    outputMemAddr <= _T_106;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (inputBlockReadable) begin
      if (isInit) begin
        if (_T_120) begin
          outputLenAddr <= _T_122;
        end else begin
          if (_T_114) begin
            outputLenAddr <= _T_118;
          end else begin
            if (_T_108) begin
              outputLenAddr <= _T_112;
            end else begin
              if (_T_104) begin
                outputLenAddr <= _T_106;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      inputAddressAccepted <= 1'h0;
    end else begin
      if (inputBlockReadable) begin
        if (_T_124) begin
          inputAddressAccepted <= 1'h0;
        end else begin
          if (_T_50) begin
            inputAddressAccepted <= 1'h1;
          end
        end
      end else begin
        if (_T_50) begin
          inputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_199) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_165) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_199) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_50 & _T_53) begin
          $fwrite(32'h80000002,"input address 0x%h accepted for core 1\n",io_inputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_165 & _T_53) begin
          $fwrite(32'h80000002,"output address 0x%h accepted for core 1\n",io_outputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module StreamingWrapper(
  input          clock,
  input          reset,
  output [63:0]  io_inputMemAddrs_0,
  output [63:0]  io_inputMemAddrs_1,
  output         io_inputMemAddrValids_0,
  output         io_inputMemAddrValids_1,
  input          io_inputMemAddrReadys_0,
  input          io_inputMemAddrReadys_1,
  input  [511:0] io_inputMemBlocks_0,
  input  [511:0] io_inputMemBlocks_1,
  input          io_inputMemBlockValids_0,
  input          io_inputMemBlockValids_1,
  output         io_inputMemBlockReadys_0,
  output         io_inputMemBlockReadys_1,
  output [63:0]  io_outputMemAddrs_0,
  output [63:0]  io_outputMemAddrs_1,
  output         io_outputMemAddrValids_0,
  output         io_outputMemAddrValids_1,
  input          io_outputMemAddrReadys_0,
  input          io_outputMemAddrReadys_1,
  output [511:0] io_outputMemBlocks_0,
  output [511:0] io_outputMemBlocks_1,
  output         io_outputMemBlockValids_0,
  output         io_outputMemBlockValids_1,
  input          io_outputMemBlockReadys_0,
  input          io_outputMemBlockReadys_1,
  output         io_finished
);
  wire  StreamingCore_clock;
  wire  StreamingCore_reset;
  wire [63:0] StreamingCore_io_inputMemAddr;
  wire  StreamingCore_io_inputMemAddrValid;
  wire  StreamingCore_io_inputMemAddrReady;
  wire [15:0] StreamingCore_io_inputMemBlock;
  wire [4:0] StreamingCore_io_inputMemIdx;
  wire  StreamingCore_io_inputMemBlockValid;
  wire  StreamingCore_io_inputMemBlockReady;
  wire [63:0] StreamingCore_io_outputMemAddr;
  wire  StreamingCore_io_outputMemAddrValid;
  wire  StreamingCore_io_outputMemAddrReady;
  wire [15:0] StreamingCore_io_outputMemBlock;
  wire [4:0] StreamingCore_io_outputMemIdx;
  wire  StreamingCore_io_outputMemBlockValid;
  wire  StreamingCore_io_outputMemBlockReady;
  wire  StreamingCore_io_inputFinished;
  wire  StreamingCore_io_outputFinished;
  wire  StreamingCore_1_clock;
  wire  StreamingCore_1_reset;
  wire [63:0] StreamingCore_1_io_inputMemAddr;
  wire  StreamingCore_1_io_inputMemAddrValid;
  wire  StreamingCore_1_io_inputMemAddrReady;
  wire [15:0] StreamingCore_1_io_inputMemBlock;
  wire [4:0] StreamingCore_1_io_inputMemIdx;
  wire  StreamingCore_1_io_inputMemBlockValid;
  wire  StreamingCore_1_io_inputMemBlockReady;
  wire [63:0] StreamingCore_1_io_outputMemAddr;
  wire  StreamingCore_1_io_outputMemAddrValid;
  wire  StreamingCore_1_io_outputMemAddrReady;
  wire [15:0] StreamingCore_1_io_outputMemBlock;
  wire [4:0] StreamingCore_1_io_outputMemIdx;
  wire  StreamingCore_1_io_outputMemBlockValid;
  wire  StreamingCore_1_io_outputMemBlockReady;
  wire  StreamingCore_1_io_inputFinished;
  wire  StreamingCore_1_io_outputFinished;
  wire [63:0] cores_0_inputMemAddr;
  wire  cores_0_inputMemAddrValid;
  wire  cores_0_inputMemAddrReady;
  wire [15:0] cores_0_inputMemBlock;
  wire [4:0] cores_0_inputMemIdx;
  wire  cores_0_inputMemBlockValid;
  wire  cores_0_inputMemBlockReady;
  wire [63:0] cores_0_outputMemAddr;
  wire  cores_0_outputMemAddrValid;
  wire  cores_0_outputMemAddrReady;
  wire [15:0] cores_0_outputMemBlock;
  wire [4:0] cores_0_outputMemIdx;
  wire  cores_0_outputMemBlockValid;
  wire  cores_0_outputMemBlockReady;
  wire  cores_0_inputFinished;
  wire  cores_0_outputFinished;
  wire [63:0] cores_1_inputMemAddr;
  wire  cores_1_inputMemAddrValid;
  wire  cores_1_inputMemAddrReady;
  wire [15:0] cores_1_inputMemBlock;
  wire [4:0] cores_1_inputMemIdx;
  wire  cores_1_inputMemBlockValid;
  wire  cores_1_inputMemBlockReady;
  wire [63:0] cores_1_outputMemAddr;
  wire  cores_1_outputMemAddrValid;
  wire  cores_1_outputMemAddrReady;
  wire [15:0] cores_1_outputMemBlock;
  wire [4:0] cores_1_outputMemIdx;
  wire  cores_1_outputMemBlockValid;
  wire  cores_1_outputMemBlockReady;
  wire  cores_1_inputFinished;
  wire  cores_1_outputFinished;
  reg  _T_239;
  reg [31:0] _RAND_0;
  reg  _T_242;
  reg [31:0] _RAND_1;
  reg  _T_245;
  reg [31:0] _RAND_2;
  reg  _T_248;
  reg [31:0] _RAND_3;
  reg [15:0] _T_252_0;
  reg [31:0] _RAND_4;
  reg [15:0] _T_252_1;
  reg [31:0] _RAND_5;
  reg [15:0] _T_252_2;
  reg [31:0] _RAND_6;
  reg [15:0] _T_252_3;
  reg [31:0] _RAND_7;
  reg [15:0] _T_252_4;
  reg [31:0] _RAND_8;
  reg [15:0] _T_252_5;
  reg [31:0] _RAND_9;
  reg [15:0] _T_252_6;
  reg [31:0] _RAND_10;
  reg [15:0] _T_252_7;
  reg [31:0] _RAND_11;
  reg [15:0] _T_252_8;
  reg [31:0] _RAND_12;
  reg [15:0] _T_252_9;
  reg [31:0] _RAND_13;
  reg [15:0] _T_252_10;
  reg [31:0] _RAND_14;
  reg [15:0] _T_252_11;
  reg [31:0] _RAND_15;
  reg [15:0] _T_252_12;
  reg [31:0] _RAND_16;
  reg [15:0] _T_252_13;
  reg [31:0] _RAND_17;
  reg [15:0] _T_252_14;
  reg [31:0] _RAND_18;
  reg [15:0] _T_252_15;
  reg [31:0] _RAND_19;
  reg [15:0] _T_252_16;
  reg [31:0] _RAND_20;
  reg [15:0] _T_252_17;
  reg [31:0] _RAND_21;
  reg [15:0] _T_252_18;
  reg [31:0] _RAND_22;
  reg [15:0] _T_252_19;
  reg [31:0] _RAND_23;
  reg [15:0] _T_252_20;
  reg [31:0] _RAND_24;
  reg [15:0] _T_252_21;
  reg [31:0] _RAND_25;
  reg [15:0] _T_252_22;
  reg [31:0] _RAND_26;
  reg [15:0] _T_252_23;
  reg [31:0] _RAND_27;
  reg [15:0] _T_252_24;
  reg [31:0] _RAND_28;
  reg [15:0] _T_252_25;
  reg [31:0] _RAND_29;
  reg [15:0] _T_252_26;
  reg [31:0] _RAND_30;
  reg [15:0] _T_252_27;
  reg [31:0] _RAND_31;
  reg [15:0] _T_252_28;
  reg [31:0] _RAND_32;
  reg [15:0] _T_252_29;
  reg [31:0] _RAND_33;
  reg [15:0] _T_252_30;
  reg [31:0] _RAND_34;
  reg [15:0] _T_252_31;
  reg [31:0] _RAND_35;
  reg [4:0] _T_289;
  reg [31:0] _RAND_36;
  reg  _T_292;
  reg [31:0] _RAND_37;
  wire  _T_293;
  wire [15:0] _T_294;
  wire [15:0] _T_295;
  wire [15:0] _T_296;
  wire [15:0] _T_297;
  wire [15:0] _T_298;
  wire [15:0] _T_299;
  wire [15:0] _T_300;
  wire [15:0] _T_301;
  wire [15:0] _T_302;
  wire [15:0] _T_303;
  wire [15:0] _T_304;
  wire [15:0] _T_305;
  wire [15:0] _T_306;
  wire [15:0] _T_307;
  wire [15:0] _T_308;
  wire [15:0] _T_309;
  wire [15:0] _T_310;
  wire [15:0] _T_311;
  wire [15:0] _T_312;
  wire [15:0] _T_313;
  wire [15:0] _T_314;
  wire [15:0] _T_315;
  wire [15:0] _T_316;
  wire [15:0] _T_317;
  wire [15:0] _T_318;
  wire [15:0] _T_319;
  wire [15:0] _T_320;
  wire [15:0] _T_321;
  wire [15:0] _T_322;
  wire [15:0] _T_323;
  wire [15:0] _T_324;
  wire [15:0] _T_325;
  wire  _T_329;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  wire [15:0] _GEN_32;
  wire [15:0] _GEN_33;
  wire [15:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire [15:0] _GEN_36;
  wire [15:0] _GEN_37;
  wire [15:0] _GEN_38;
  wire [15:0] _GEN_39;
  wire [15:0] _GEN_40;
  wire [15:0] _GEN_41;
  wire [15:0] _GEN_42;
  wire [15:0] _GEN_43;
  wire [15:0] _GEN_44;
  wire [15:0] _GEN_45;
  wire [15:0] _GEN_46;
  wire [15:0] _GEN_47;
  wire [15:0] _GEN_48;
  wire [15:0] _GEN_49;
  wire [15:0] _GEN_50;
  wire [15:0] _GEN_51;
  wire [15:0] _GEN_52;
  wire [15:0] _GEN_53;
  wire [15:0] _GEN_54;
  wire [15:0] _GEN_55;
  wire [15:0] _GEN_56;
  wire [15:0] _GEN_57;
  wire  _GEN_58;
  wire  _T_331;
  wire [5:0] _T_335;
  wire [4:0] _T_336;
  wire  _GEN_59;
  wire [4:0] _GEN_60;
  wire  _GEN_61;
  wire [4:0] _GEN_62;
  wire [63:0] _GEN_0_inputMemAddr;
  wire [63:0] _GEN_63;
  wire  _GEN_64;
  wire  _GEN_69;
  wire  _GEN_77;
  wire  _GEN_1_inputMemAddrValid;
  wire  _GEN_2_inputMemBlockReady;
  wire  _T_437;
  wire  _T_439;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_79;
  wire [15:0] _GEN_80;
  wire [15:0] _GEN_81;
  wire [15:0] _GEN_82;
  wire [15:0] _GEN_83;
  wire [15:0] _GEN_84;
  wire [15:0] _GEN_85;
  wire [15:0] _GEN_86;
  wire [15:0] _GEN_87;
  wire [15:0] _GEN_88;
  wire [15:0] _GEN_89;
  wire [15:0] _GEN_90;
  wire [15:0] _GEN_91;
  wire [15:0] _GEN_92;
  wire [15:0] _GEN_93;
  wire [15:0] _GEN_94;
  wire [15:0] _GEN_95;
  wire [15:0] _GEN_96;
  wire [15:0] _GEN_97;
  wire [15:0] _GEN_98;
  wire [15:0] _GEN_99;
  wire [15:0] _GEN_100;
  wire [15:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire [15:0] _GEN_103;
  wire [15:0] _GEN_104;
  wire [15:0] _GEN_105;
  wire [15:0] _GEN_106;
  wire [15:0] _GEN_107;
  wire [15:0] _GEN_108;
  wire [15:0] _GEN_109;
  wire  _T_444;
  wire  _GEN_4_inputFinished;
  wire  _T_480;
  wire [1:0] _T_485;
  wire  _T_486;
  wire  _T_487;
  wire  _GEN_110;
  reg [15:0] _T_491_0;
  reg [31:0] _RAND_38;
  reg [15:0] _T_491_1;
  reg [31:0] _RAND_39;
  reg [15:0] _T_491_2;
  reg [31:0] _RAND_40;
  reg [15:0] _T_491_3;
  reg [31:0] _RAND_41;
  reg [15:0] _T_491_4;
  reg [31:0] _RAND_42;
  reg [15:0] _T_491_5;
  reg [31:0] _RAND_43;
  reg [15:0] _T_491_6;
  reg [31:0] _RAND_44;
  reg [15:0] _T_491_7;
  reg [31:0] _RAND_45;
  reg [15:0] _T_491_8;
  reg [31:0] _RAND_46;
  reg [15:0] _T_491_9;
  reg [31:0] _RAND_47;
  reg [15:0] _T_491_10;
  reg [31:0] _RAND_48;
  reg [15:0] _T_491_11;
  reg [31:0] _RAND_49;
  reg [15:0] _T_491_12;
  reg [31:0] _RAND_50;
  reg [15:0] _T_491_13;
  reg [31:0] _RAND_51;
  reg [15:0] _T_491_14;
  reg [31:0] _RAND_52;
  reg [15:0] _T_491_15;
  reg [31:0] _RAND_53;
  reg [15:0] _T_491_16;
  reg [31:0] _RAND_54;
  reg [15:0] _T_491_17;
  reg [31:0] _RAND_55;
  reg [15:0] _T_491_18;
  reg [31:0] _RAND_56;
  reg [15:0] _T_491_19;
  reg [31:0] _RAND_57;
  reg [15:0] _T_491_20;
  reg [31:0] _RAND_58;
  reg [15:0] _T_491_21;
  reg [31:0] _RAND_59;
  reg [15:0] _T_491_22;
  reg [31:0] _RAND_60;
  reg [15:0] _T_491_23;
  reg [31:0] _RAND_61;
  reg [15:0] _T_491_24;
  reg [31:0] _RAND_62;
  reg [15:0] _T_491_25;
  reg [31:0] _RAND_63;
  reg [15:0] _T_491_26;
  reg [31:0] _RAND_64;
  reg [15:0] _T_491_27;
  reg [31:0] _RAND_65;
  reg [15:0] _T_491_28;
  reg [31:0] _RAND_66;
  reg [15:0] _T_491_29;
  reg [31:0] _RAND_67;
  reg [15:0] _T_491_30;
  reg [31:0] _RAND_68;
  reg [15:0] _T_491_31;
  reg [31:0] _RAND_69;
  reg [4:0] _T_528;
  reg [31:0] _RAND_70;
  reg  _T_531;
  reg [31:0] _RAND_71;
  wire  _T_532;
  wire [15:0] _T_533;
  wire [15:0] _T_534;
  wire [15:0] _T_535;
  wire [15:0] _T_536;
  wire [15:0] _T_537;
  wire [15:0] _T_538;
  wire [15:0] _T_539;
  wire [15:0] _T_540;
  wire [15:0] _T_541;
  wire [15:0] _T_542;
  wire [15:0] _T_543;
  wire [15:0] _T_544;
  wire [15:0] _T_545;
  wire [15:0] _T_546;
  wire [15:0] _T_547;
  wire [15:0] _T_548;
  wire [15:0] _T_549;
  wire [15:0] _T_550;
  wire [15:0] _T_551;
  wire [15:0] _T_552;
  wire [15:0] _T_553;
  wire [15:0] _T_554;
  wire [15:0] _T_555;
  wire [15:0] _T_556;
  wire [15:0] _T_557;
  wire [15:0] _T_558;
  wire [15:0] _T_559;
  wire [15:0] _T_560;
  wire [15:0] _T_561;
  wire [15:0] _T_562;
  wire [15:0] _T_563;
  wire [15:0] _T_564;
  wire [15:0] _GEN_111;
  wire [15:0] _GEN_112;
  wire [15:0] _GEN_113;
  wire [15:0] _GEN_114;
  wire [15:0] _GEN_115;
  wire [15:0] _GEN_116;
  wire [15:0] _GEN_117;
  wire [15:0] _GEN_118;
  wire [15:0] _GEN_119;
  wire [15:0] _GEN_120;
  wire [15:0] _GEN_121;
  wire [15:0] _GEN_122;
  wire [15:0] _GEN_123;
  wire [15:0] _GEN_124;
  wire [15:0] _GEN_125;
  wire [15:0] _GEN_126;
  wire [15:0] _GEN_127;
  wire [15:0] _GEN_128;
  wire [15:0] _GEN_129;
  wire [15:0] _GEN_130;
  wire [15:0] _GEN_131;
  wire [15:0] _GEN_132;
  wire [15:0] _GEN_133;
  wire [15:0] _GEN_134;
  wire [15:0] _GEN_135;
  wire [15:0] _GEN_136;
  wire [15:0] _GEN_137;
  wire [15:0] _GEN_138;
  wire [15:0] _GEN_139;
  wire [15:0] _GEN_140;
  wire [15:0] _GEN_141;
  wire [15:0] _GEN_142;
  wire  _GEN_143;
  wire  _T_570;
  wire [5:0] _T_574;
  wire [4:0] _T_575;
  wire  _GEN_144;
  wire [4:0] _GEN_145;
  wire  _GEN_146;
  wire [4:0] _GEN_147;
  wire [63:0] _GEN_5_inputMemAddr;
  wire [63:0] _GEN_148;
  wire  _GEN_149;
  wire  _GEN_154;
  wire  _GEN_162;
  wire  _GEN_6_inputMemAddrValid;
  wire  _GEN_7_inputMemBlockReady;
  wire  _T_678;
  wire [15:0] _GEN_8;
  wire [15:0] _GEN_164;
  wire [15:0] _GEN_165;
  wire [15:0] _GEN_166;
  wire [15:0] _GEN_167;
  wire [15:0] _GEN_168;
  wire [15:0] _GEN_169;
  wire [15:0] _GEN_170;
  wire [15:0] _GEN_171;
  wire [15:0] _GEN_172;
  wire [15:0] _GEN_173;
  wire [15:0] _GEN_174;
  wire [15:0] _GEN_175;
  wire [15:0] _GEN_176;
  wire [15:0] _GEN_177;
  wire [15:0] _GEN_178;
  wire [15:0] _GEN_179;
  wire [15:0] _GEN_180;
  wire [15:0] _GEN_181;
  wire [15:0] _GEN_182;
  wire [15:0] _GEN_183;
  wire [15:0] _GEN_184;
  wire [15:0] _GEN_185;
  wire [15:0] _GEN_186;
  wire [15:0] _GEN_187;
  wire [15:0] _GEN_188;
  wire [15:0] _GEN_189;
  wire [15:0] _GEN_190;
  wire [15:0] _GEN_191;
  wire [15:0] _GEN_192;
  wire [15:0] _GEN_193;
  wire [15:0] _GEN_194;
  wire  _T_683;
  wire  _GEN_9_inputFinished;
  wire  _T_719;
  wire [1:0] _T_724;
  wire  _T_725;
  wire  _T_726;
  wire  _GEN_195;
  reg [15:0] _T_730_0;
  reg [31:0] _RAND_72;
  reg [15:0] _T_730_1;
  reg [31:0] _RAND_73;
  reg [15:0] _T_730_2;
  reg [31:0] _RAND_74;
  reg [15:0] _T_730_3;
  reg [31:0] _RAND_75;
  reg [15:0] _T_730_4;
  reg [31:0] _RAND_76;
  reg [15:0] _T_730_5;
  reg [31:0] _RAND_77;
  reg [15:0] _T_730_6;
  reg [31:0] _RAND_78;
  reg [15:0] _T_730_7;
  reg [31:0] _RAND_79;
  reg [15:0] _T_730_8;
  reg [31:0] _RAND_80;
  reg [15:0] _T_730_9;
  reg [31:0] _RAND_81;
  reg [15:0] _T_730_10;
  reg [31:0] _RAND_82;
  reg [15:0] _T_730_11;
  reg [31:0] _RAND_83;
  reg [15:0] _T_730_12;
  reg [31:0] _RAND_84;
  reg [15:0] _T_730_13;
  reg [31:0] _RAND_85;
  reg [15:0] _T_730_14;
  reg [31:0] _RAND_86;
  reg [15:0] _T_730_15;
  reg [31:0] _RAND_87;
  reg [15:0] _T_730_16;
  reg [31:0] _RAND_88;
  reg [15:0] _T_730_17;
  reg [31:0] _RAND_89;
  reg [15:0] _T_730_18;
  reg [31:0] _RAND_90;
  reg [15:0] _T_730_19;
  reg [31:0] _RAND_91;
  reg [15:0] _T_730_20;
  reg [31:0] _RAND_92;
  reg [15:0] _T_730_21;
  reg [31:0] _RAND_93;
  reg [15:0] _T_730_22;
  reg [31:0] _RAND_94;
  reg [15:0] _T_730_23;
  reg [31:0] _RAND_95;
  reg [15:0] _T_730_24;
  reg [31:0] _RAND_96;
  reg [15:0] _T_730_25;
  reg [31:0] _RAND_97;
  reg [15:0] _T_730_26;
  reg [31:0] _RAND_98;
  reg [15:0] _T_730_27;
  reg [31:0] _RAND_99;
  reg [15:0] _T_730_28;
  reg [31:0] _RAND_100;
  reg [15:0] _T_730_29;
  reg [31:0] _RAND_101;
  reg [15:0] _T_730_30;
  reg [31:0] _RAND_102;
  reg [15:0] _T_730_31;
  reg [31:0] _RAND_103;
  reg  _T_767;
  reg [31:0] _RAND_104;
  wire [4:0] _GEN_10_outputMemIdx;
  wire [63:0] _GEN_203;
  wire  _GEN_204;
  wire [15:0] _GEN_206;
  wire [4:0] _GEN_207;
  wire  _GEN_208;
  wire  _GEN_211;
  wire  _T_835;
  wire  _GEN_11_outputMemBlockValid;
  wire  _T_836;
  wire  _GEN_212;
  wire  _T_839;
  wire [4:0] _GEN_12_outputMemIdx;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_213;
  wire [15:0] _GEN_214;
  wire [15:0] _GEN_215;
  wire [15:0] _GEN_216;
  wire [15:0] _GEN_217;
  wire [15:0] _GEN_218;
  wire [15:0] _GEN_219;
  wire [15:0] _GEN_220;
  wire [15:0] _GEN_221;
  wire [15:0] _GEN_222;
  wire [15:0] _GEN_223;
  wire [15:0] _GEN_224;
  wire [15:0] _GEN_225;
  wire [15:0] _GEN_226;
  wire [15:0] _GEN_227;
  wire [15:0] _GEN_228;
  wire [15:0] _GEN_229;
  wire [15:0] _GEN_230;
  wire [15:0] _GEN_231;
  wire [15:0] _GEN_232;
  wire [15:0] _GEN_233;
  wire [15:0] _GEN_234;
  wire [15:0] _GEN_235;
  wire [15:0] _GEN_236;
  wire [15:0] _GEN_237;
  wire [15:0] _GEN_238;
  wire [15:0] _GEN_239;
  wire [15:0] _GEN_240;
  wire [15:0] _GEN_241;
  wire [15:0] _GEN_242;
  wire [15:0] _GEN_243;
  wire [15:0] _GEN_244;
  wire [15:0] _GEN_14_outputMemBlock;
  wire [15:0] _GEN_245;
  wire [15:0] _GEN_246;
  wire [15:0] _GEN_247;
  wire [15:0] _GEN_248;
  wire [15:0] _GEN_249;
  wire [15:0] _GEN_250;
  wire [15:0] _GEN_251;
  wire [15:0] _GEN_252;
  wire [15:0] _GEN_253;
  wire [15:0] _GEN_254;
  wire [15:0] _GEN_255;
  wire [15:0] _GEN_256;
  wire [15:0] _GEN_257;
  wire [15:0] _GEN_258;
  wire [15:0] _GEN_259;
  wire [15:0] _GEN_260;
  wire [15:0] _GEN_261;
  wire [15:0] _GEN_262;
  wire [15:0] _GEN_263;
  wire [15:0] _GEN_264;
  wire [15:0] _GEN_265;
  wire [15:0] _GEN_266;
  wire [15:0] _GEN_267;
  wire [15:0] _GEN_268;
  wire [15:0] _GEN_269;
  wire [15:0] _GEN_270;
  wire [15:0] _GEN_271;
  wire [15:0] _GEN_272;
  wire [15:0] _GEN_273;
  wire [15:0] _GEN_274;
  wire [15:0] _GEN_275;
  wire [15:0] _GEN_276;
  wire [63:0] _GEN_15_outputMemAddr;
  wire  _GEN_16_outputMemAddrValid;
  wire [31:0] _T_973;
  wire [31:0] _T_974;
  wire [63:0] _T_975;
  wire [31:0] _T_976;
  wire [31:0] _T_977;
  wire [63:0] _T_978;
  wire [127:0] _T_979;
  wire [31:0] _T_980;
  wire [31:0] _T_981;
  wire [63:0] _T_982;
  wire [31:0] _T_983;
  wire [31:0] _T_984;
  wire [63:0] _T_985;
  wire [127:0] _T_986;
  wire [255:0] _T_987;
  wire [31:0] _T_988;
  wire [31:0] _T_989;
  wire [63:0] _T_990;
  wire [31:0] _T_991;
  wire [31:0] _T_992;
  wire [63:0] _T_993;
  wire [127:0] _T_994;
  wire [31:0] _T_995;
  wire [31:0] _T_996;
  wire [63:0] _T_997;
  wire [31:0] _T_998;
  wire [31:0] _T_999;
  wire [63:0] _T_1000;
  wire [127:0] _T_1001;
  wire [255:0] _T_1002;
  wire [511:0] _T_1003;
  wire  _T_1005;
  wire  _T_1007;
  wire  _T_1010;
  wire  _T_1012;
  wire  _T_1013;
  wire  _GEN_17_outputFinished;
  wire  _T_1051;
  wire [1:0] _T_1056;
  wire  _T_1057;
  wire  _T_1058;
  wire  _GEN_277;
  wire  _GEN_278;
  reg [15:0] _T_1063_0;
  reg [31:0] _RAND_105;
  reg [15:0] _T_1063_1;
  reg [31:0] _RAND_106;
  reg [15:0] _T_1063_2;
  reg [31:0] _RAND_107;
  reg [15:0] _T_1063_3;
  reg [31:0] _RAND_108;
  reg [15:0] _T_1063_4;
  reg [31:0] _RAND_109;
  reg [15:0] _T_1063_5;
  reg [31:0] _RAND_110;
  reg [15:0] _T_1063_6;
  reg [31:0] _RAND_111;
  reg [15:0] _T_1063_7;
  reg [31:0] _RAND_112;
  reg [15:0] _T_1063_8;
  reg [31:0] _RAND_113;
  reg [15:0] _T_1063_9;
  reg [31:0] _RAND_114;
  reg [15:0] _T_1063_10;
  reg [31:0] _RAND_115;
  reg [15:0] _T_1063_11;
  reg [31:0] _RAND_116;
  reg [15:0] _T_1063_12;
  reg [31:0] _RAND_117;
  reg [15:0] _T_1063_13;
  reg [31:0] _RAND_118;
  reg [15:0] _T_1063_14;
  reg [31:0] _RAND_119;
  reg [15:0] _T_1063_15;
  reg [31:0] _RAND_120;
  reg [15:0] _T_1063_16;
  reg [31:0] _RAND_121;
  reg [15:0] _T_1063_17;
  reg [31:0] _RAND_122;
  reg [15:0] _T_1063_18;
  reg [31:0] _RAND_123;
  reg [15:0] _T_1063_19;
  reg [31:0] _RAND_124;
  reg [15:0] _T_1063_20;
  reg [31:0] _RAND_125;
  reg [15:0] _T_1063_21;
  reg [31:0] _RAND_126;
  reg [15:0] _T_1063_22;
  reg [31:0] _RAND_127;
  reg [15:0] _T_1063_23;
  reg [31:0] _RAND_128;
  reg [15:0] _T_1063_24;
  reg [31:0] _RAND_129;
  reg [15:0] _T_1063_25;
  reg [31:0] _RAND_130;
  reg [15:0] _T_1063_26;
  reg [31:0] _RAND_131;
  reg [15:0] _T_1063_27;
  reg [31:0] _RAND_132;
  reg [15:0] _T_1063_28;
  reg [31:0] _RAND_133;
  reg [15:0] _T_1063_29;
  reg [31:0] _RAND_134;
  reg [15:0] _T_1063_30;
  reg [31:0] _RAND_135;
  reg [15:0] _T_1063_31;
  reg [31:0] _RAND_136;
  reg  _T_1100;
  reg [31:0] _RAND_137;
  wire [4:0] _GEN_18_outputMemIdx;
  wire [63:0] _GEN_286;
  wire  _GEN_287;
  wire [15:0] _GEN_289;
  wire [4:0] _GEN_290;
  wire  _GEN_291;
  wire  _GEN_294;
  wire  _T_1168;
  wire  _GEN_19_outputMemBlockValid;
  wire  _T_1169;
  wire  _GEN_295;
  wire  _T_1172;
  wire [4:0] _GEN_20_outputMemIdx;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_296;
  wire [15:0] _GEN_297;
  wire [15:0] _GEN_298;
  wire [15:0] _GEN_299;
  wire [15:0] _GEN_300;
  wire [15:0] _GEN_301;
  wire [15:0] _GEN_302;
  wire [15:0] _GEN_303;
  wire [15:0] _GEN_304;
  wire [15:0] _GEN_305;
  wire [15:0] _GEN_306;
  wire [15:0] _GEN_307;
  wire [15:0] _GEN_308;
  wire [15:0] _GEN_309;
  wire [15:0] _GEN_310;
  wire [15:0] _GEN_311;
  wire [15:0] _GEN_312;
  wire [15:0] _GEN_313;
  wire [15:0] _GEN_314;
  wire [15:0] _GEN_315;
  wire [15:0] _GEN_316;
  wire [15:0] _GEN_317;
  wire [15:0] _GEN_318;
  wire [15:0] _GEN_319;
  wire [15:0] _GEN_320;
  wire [15:0] _GEN_321;
  wire [15:0] _GEN_322;
  wire [15:0] _GEN_323;
  wire [15:0] _GEN_324;
  wire [15:0] _GEN_325;
  wire [15:0] _GEN_326;
  wire [15:0] _GEN_327;
  wire [15:0] _GEN_22_outputMemBlock;
  wire [15:0] _GEN_328;
  wire [15:0] _GEN_329;
  wire [15:0] _GEN_330;
  wire [15:0] _GEN_331;
  wire [15:0] _GEN_332;
  wire [15:0] _GEN_333;
  wire [15:0] _GEN_334;
  wire [15:0] _GEN_335;
  wire [15:0] _GEN_336;
  wire [15:0] _GEN_337;
  wire [15:0] _GEN_338;
  wire [15:0] _GEN_339;
  wire [15:0] _GEN_340;
  wire [15:0] _GEN_341;
  wire [15:0] _GEN_342;
  wire [15:0] _GEN_343;
  wire [15:0] _GEN_344;
  wire [15:0] _GEN_345;
  wire [15:0] _GEN_346;
  wire [15:0] _GEN_347;
  wire [15:0] _GEN_348;
  wire [15:0] _GEN_349;
  wire [15:0] _GEN_350;
  wire [15:0] _GEN_351;
  wire [15:0] _GEN_352;
  wire [15:0] _GEN_353;
  wire [15:0] _GEN_354;
  wire [15:0] _GEN_355;
  wire [15:0] _GEN_356;
  wire [15:0] _GEN_357;
  wire [15:0] _GEN_358;
  wire [15:0] _GEN_359;
  wire [63:0] _GEN_23_outputMemAddr;
  wire  _GEN_24_outputMemAddrValid;
  wire [31:0] _T_1306;
  wire [31:0] _T_1307;
  wire [63:0] _T_1308;
  wire [31:0] _T_1309;
  wire [31:0] _T_1310;
  wire [63:0] _T_1311;
  wire [127:0] _T_1312;
  wire [31:0] _T_1313;
  wire [31:0] _T_1314;
  wire [63:0] _T_1315;
  wire [31:0] _T_1316;
  wire [31:0] _T_1317;
  wire [63:0] _T_1318;
  wire [127:0] _T_1319;
  wire [255:0] _T_1320;
  wire [31:0] _T_1321;
  wire [31:0] _T_1322;
  wire [63:0] _T_1323;
  wire [31:0] _T_1324;
  wire [31:0] _T_1325;
  wire [63:0] _T_1326;
  wire [127:0] _T_1327;
  wire [31:0] _T_1328;
  wire [31:0] _T_1329;
  wire [63:0] _T_1330;
  wire [31:0] _T_1331;
  wire [31:0] _T_1332;
  wire [63:0] _T_1333;
  wire [127:0] _T_1334;
  wire [255:0] _T_1335;
  wire [511:0] _T_1336;
  wire  _T_1340;
  wire  _T_1343;
  wire  _T_1345;
  wire  _T_1346;
  wire  _GEN_25_outputFinished;
  wire  _T_1384;
  wire [1:0] _T_1389;
  wire  _T_1390;
  wire  _T_1391;
  wire  _GEN_360;
  wire  _GEN_361;
  wire  cumFinished;
  StreamingCore StreamingCore (
    .clock(StreamingCore_clock),
    .reset(StreamingCore_reset),
    .io_inputMemAddr(StreamingCore_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_io_inputMemAddrValid),
    .io_inputMemAddrReady(StreamingCore_io_inputMemAddrReady),
    .io_inputMemBlock(StreamingCore_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_io_outputMemBlockReady),
    .io_inputFinished(StreamingCore_io_inputFinished),
    .io_outputFinished(StreamingCore_io_outputFinished)
  );
  StreamingCore_1 StreamingCore_1 (
    .clock(StreamingCore_1_clock),
    .reset(StreamingCore_1_reset),
    .io_inputMemAddr(StreamingCore_1_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_1_io_inputMemAddrValid),
    .io_inputMemAddrReady(StreamingCore_1_io_inputMemAddrReady),
    .io_inputMemBlock(StreamingCore_1_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_1_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_1_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_1_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_1_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_1_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_1_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_1_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_1_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_1_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_1_io_outputMemBlockReady),
    .io_inputFinished(StreamingCore_1_io_inputFinished),
    .io_outputFinished(StreamingCore_1_io_outputFinished)
  );
  assign _T_293 = io_inputMemBlockReadys_0 & io_inputMemBlockValids_0;
  assign _T_294 = io_inputMemBlocks_0[15:0];
  assign _T_295 = io_inputMemBlocks_0[31:16];
  assign _T_296 = io_inputMemBlocks_0[47:32];
  assign _T_297 = io_inputMemBlocks_0[63:48];
  assign _T_298 = io_inputMemBlocks_0[79:64];
  assign _T_299 = io_inputMemBlocks_0[95:80];
  assign _T_300 = io_inputMemBlocks_0[111:96];
  assign _T_301 = io_inputMemBlocks_0[127:112];
  assign _T_302 = io_inputMemBlocks_0[143:128];
  assign _T_303 = io_inputMemBlocks_0[159:144];
  assign _T_304 = io_inputMemBlocks_0[175:160];
  assign _T_305 = io_inputMemBlocks_0[191:176];
  assign _T_306 = io_inputMemBlocks_0[207:192];
  assign _T_307 = io_inputMemBlocks_0[223:208];
  assign _T_308 = io_inputMemBlocks_0[239:224];
  assign _T_309 = io_inputMemBlocks_0[255:240];
  assign _T_310 = io_inputMemBlocks_0[271:256];
  assign _T_311 = io_inputMemBlocks_0[287:272];
  assign _T_312 = io_inputMemBlocks_0[303:288];
  assign _T_313 = io_inputMemBlocks_0[319:304];
  assign _T_314 = io_inputMemBlocks_0[335:320];
  assign _T_315 = io_inputMemBlocks_0[351:336];
  assign _T_316 = io_inputMemBlocks_0[367:352];
  assign _T_317 = io_inputMemBlocks_0[383:368];
  assign _T_318 = io_inputMemBlocks_0[399:384];
  assign _T_319 = io_inputMemBlocks_0[415:400];
  assign _T_320 = io_inputMemBlocks_0[431:416];
  assign _T_321 = io_inputMemBlocks_0[447:432];
  assign _T_322 = io_inputMemBlocks_0[463:448];
  assign _T_323 = io_inputMemBlocks_0[479:464];
  assign _T_324 = io_inputMemBlocks_0[495:480];
  assign _T_325 = io_inputMemBlocks_0[511:496];
  assign _T_329 = reset == 1'h0;
  assign _GEN_26 = _T_293 ? _T_294 : _T_252_0;
  assign _GEN_27 = _T_293 ? _T_295 : _T_252_1;
  assign _GEN_28 = _T_293 ? _T_296 : _T_252_2;
  assign _GEN_29 = _T_293 ? _T_297 : _T_252_3;
  assign _GEN_30 = _T_293 ? _T_298 : _T_252_4;
  assign _GEN_31 = _T_293 ? _T_299 : _T_252_5;
  assign _GEN_32 = _T_293 ? _T_300 : _T_252_6;
  assign _GEN_33 = _T_293 ? _T_301 : _T_252_7;
  assign _GEN_34 = _T_293 ? _T_302 : _T_252_8;
  assign _GEN_35 = _T_293 ? _T_303 : _T_252_9;
  assign _GEN_36 = _T_293 ? _T_304 : _T_252_10;
  assign _GEN_37 = _T_293 ? _T_305 : _T_252_11;
  assign _GEN_38 = _T_293 ? _T_306 : _T_252_12;
  assign _GEN_39 = _T_293 ? _T_307 : _T_252_13;
  assign _GEN_40 = _T_293 ? _T_308 : _T_252_14;
  assign _GEN_41 = _T_293 ? _T_309 : _T_252_15;
  assign _GEN_42 = _T_293 ? _T_310 : _T_252_16;
  assign _GEN_43 = _T_293 ? _T_311 : _T_252_17;
  assign _GEN_44 = _T_293 ? _T_312 : _T_252_18;
  assign _GEN_45 = _T_293 ? _T_313 : _T_252_19;
  assign _GEN_46 = _T_293 ? _T_314 : _T_252_20;
  assign _GEN_47 = _T_293 ? _T_315 : _T_252_21;
  assign _GEN_48 = _T_293 ? _T_316 : _T_252_22;
  assign _GEN_49 = _T_293 ? _T_317 : _T_252_23;
  assign _GEN_50 = _T_293 ? _T_318 : _T_252_24;
  assign _GEN_51 = _T_293 ? _T_319 : _T_252_25;
  assign _GEN_52 = _T_293 ? _T_320 : _T_252_26;
  assign _GEN_53 = _T_293 ? _T_321 : _T_252_27;
  assign _GEN_54 = _T_293 ? _T_322 : _T_252_28;
  assign _GEN_55 = _T_293 ? _T_323 : _T_252_29;
  assign _GEN_56 = _T_293 ? _T_324 : _T_252_30;
  assign _GEN_57 = _T_293 ? _T_325 : _T_252_31;
  assign _GEN_58 = _T_293 ? 1'h1 : _T_292;
  assign _T_331 = _T_289 == 5'h1f;
  assign _T_335 = _T_289 + 5'h1;
  assign _T_336 = _T_335[4:0];
  assign _GEN_59 = _T_331 ? 1'h0 : _GEN_58;
  assign _GEN_60 = _T_331 ? 5'h0 : _T_336;
  assign _GEN_61 = _T_292 ? _GEN_59 : _GEN_58;
  assign _GEN_62 = _T_292 ? _GEN_60 : _T_289;
  assign _GEN_63 = _T_239 ? cores_1_inputMemAddr : cores_0_inputMemAddr;
  assign _GEN_64 = _T_239 ? cores_1_inputMemAddrValid : cores_0_inputMemAddrValid;
  assign _GEN_69 = _T_239 ? cores_1_inputMemBlockReady : cores_0_inputMemBlockReady;
  assign _GEN_77 = _T_239 ? cores_1_inputFinished : cores_0_inputFinished;
  assign _T_437 = _T_239 == 1'h0;
  assign _T_439 = _T_437 ? io_inputMemAddrReadys_0 : 1'h0;
  assign _GEN_79 = 5'h1 == _T_289 ? _T_252_1 : _T_252_0;
  assign _GEN_80 = 5'h2 == _T_289 ? _T_252_2 : _GEN_79;
  assign _GEN_81 = 5'h3 == _T_289 ? _T_252_3 : _GEN_80;
  assign _GEN_82 = 5'h4 == _T_289 ? _T_252_4 : _GEN_81;
  assign _GEN_83 = 5'h5 == _T_289 ? _T_252_5 : _GEN_82;
  assign _GEN_84 = 5'h6 == _T_289 ? _T_252_6 : _GEN_83;
  assign _GEN_85 = 5'h7 == _T_289 ? _T_252_7 : _GEN_84;
  assign _GEN_86 = 5'h8 == _T_289 ? _T_252_8 : _GEN_85;
  assign _GEN_87 = 5'h9 == _T_289 ? _T_252_9 : _GEN_86;
  assign _GEN_88 = 5'ha == _T_289 ? _T_252_10 : _GEN_87;
  assign _GEN_89 = 5'hb == _T_289 ? _T_252_11 : _GEN_88;
  assign _GEN_90 = 5'hc == _T_289 ? _T_252_12 : _GEN_89;
  assign _GEN_91 = 5'hd == _T_289 ? _T_252_13 : _GEN_90;
  assign _GEN_92 = 5'he == _T_289 ? _T_252_14 : _GEN_91;
  assign _GEN_93 = 5'hf == _T_289 ? _T_252_15 : _GEN_92;
  assign _GEN_94 = 5'h10 == _T_289 ? _T_252_16 : _GEN_93;
  assign _GEN_95 = 5'h11 == _T_289 ? _T_252_17 : _GEN_94;
  assign _GEN_96 = 5'h12 == _T_289 ? _T_252_18 : _GEN_95;
  assign _GEN_97 = 5'h13 == _T_289 ? _T_252_19 : _GEN_96;
  assign _GEN_98 = 5'h14 == _T_289 ? _T_252_20 : _GEN_97;
  assign _GEN_99 = 5'h15 == _T_289 ? _T_252_21 : _GEN_98;
  assign _GEN_100 = 5'h16 == _T_289 ? _T_252_22 : _GEN_99;
  assign _GEN_101 = 5'h17 == _T_289 ? _T_252_23 : _GEN_100;
  assign _GEN_102 = 5'h18 == _T_289 ? _T_252_24 : _GEN_101;
  assign _GEN_103 = 5'h19 == _T_289 ? _T_252_25 : _GEN_102;
  assign _GEN_104 = 5'h1a == _T_289 ? _T_252_26 : _GEN_103;
  assign _GEN_105 = 5'h1b == _T_289 ? _T_252_27 : _GEN_104;
  assign _GEN_106 = 5'h1c == _T_289 ? _T_252_28 : _GEN_105;
  assign _GEN_107 = 5'h1d == _T_289 ? _T_252_29 : _GEN_106;
  assign _GEN_108 = 5'h1e == _T_289 ? _T_252_30 : _GEN_107;
  assign _GEN_109 = 5'h1f == _T_289 ? _T_252_31 : _GEN_108;
  assign _T_444 = _T_437 ? _T_292 : 1'h0;
  assign _T_480 = _GEN_4_inputFinished | _T_331;
  assign _T_485 = _T_239 + 1'h1;
  assign _T_486 = _T_485[0:0];
  assign _T_487 = _T_437 ? 1'h0 : _T_486;
  assign _GEN_110 = _T_480 ? _T_487 : _T_239;
  assign _T_532 = io_inputMemBlockReadys_1 & io_inputMemBlockValids_1;
  assign _T_533 = io_inputMemBlocks_1[15:0];
  assign _T_534 = io_inputMemBlocks_1[31:16];
  assign _T_535 = io_inputMemBlocks_1[47:32];
  assign _T_536 = io_inputMemBlocks_1[63:48];
  assign _T_537 = io_inputMemBlocks_1[79:64];
  assign _T_538 = io_inputMemBlocks_1[95:80];
  assign _T_539 = io_inputMemBlocks_1[111:96];
  assign _T_540 = io_inputMemBlocks_1[127:112];
  assign _T_541 = io_inputMemBlocks_1[143:128];
  assign _T_542 = io_inputMemBlocks_1[159:144];
  assign _T_543 = io_inputMemBlocks_1[175:160];
  assign _T_544 = io_inputMemBlocks_1[191:176];
  assign _T_545 = io_inputMemBlocks_1[207:192];
  assign _T_546 = io_inputMemBlocks_1[223:208];
  assign _T_547 = io_inputMemBlocks_1[239:224];
  assign _T_548 = io_inputMemBlocks_1[255:240];
  assign _T_549 = io_inputMemBlocks_1[271:256];
  assign _T_550 = io_inputMemBlocks_1[287:272];
  assign _T_551 = io_inputMemBlocks_1[303:288];
  assign _T_552 = io_inputMemBlocks_1[319:304];
  assign _T_553 = io_inputMemBlocks_1[335:320];
  assign _T_554 = io_inputMemBlocks_1[351:336];
  assign _T_555 = io_inputMemBlocks_1[367:352];
  assign _T_556 = io_inputMemBlocks_1[383:368];
  assign _T_557 = io_inputMemBlocks_1[399:384];
  assign _T_558 = io_inputMemBlocks_1[415:400];
  assign _T_559 = io_inputMemBlocks_1[431:416];
  assign _T_560 = io_inputMemBlocks_1[447:432];
  assign _T_561 = io_inputMemBlocks_1[463:448];
  assign _T_562 = io_inputMemBlocks_1[479:464];
  assign _T_563 = io_inputMemBlocks_1[495:480];
  assign _T_564 = io_inputMemBlocks_1[511:496];
  assign _GEN_111 = _T_532 ? _T_533 : _T_491_0;
  assign _GEN_112 = _T_532 ? _T_534 : _T_491_1;
  assign _GEN_113 = _T_532 ? _T_535 : _T_491_2;
  assign _GEN_114 = _T_532 ? _T_536 : _T_491_3;
  assign _GEN_115 = _T_532 ? _T_537 : _T_491_4;
  assign _GEN_116 = _T_532 ? _T_538 : _T_491_5;
  assign _GEN_117 = _T_532 ? _T_539 : _T_491_6;
  assign _GEN_118 = _T_532 ? _T_540 : _T_491_7;
  assign _GEN_119 = _T_532 ? _T_541 : _T_491_8;
  assign _GEN_120 = _T_532 ? _T_542 : _T_491_9;
  assign _GEN_121 = _T_532 ? _T_543 : _T_491_10;
  assign _GEN_122 = _T_532 ? _T_544 : _T_491_11;
  assign _GEN_123 = _T_532 ? _T_545 : _T_491_12;
  assign _GEN_124 = _T_532 ? _T_546 : _T_491_13;
  assign _GEN_125 = _T_532 ? _T_547 : _T_491_14;
  assign _GEN_126 = _T_532 ? _T_548 : _T_491_15;
  assign _GEN_127 = _T_532 ? _T_549 : _T_491_16;
  assign _GEN_128 = _T_532 ? _T_550 : _T_491_17;
  assign _GEN_129 = _T_532 ? _T_551 : _T_491_18;
  assign _GEN_130 = _T_532 ? _T_552 : _T_491_19;
  assign _GEN_131 = _T_532 ? _T_553 : _T_491_20;
  assign _GEN_132 = _T_532 ? _T_554 : _T_491_21;
  assign _GEN_133 = _T_532 ? _T_555 : _T_491_22;
  assign _GEN_134 = _T_532 ? _T_556 : _T_491_23;
  assign _GEN_135 = _T_532 ? _T_557 : _T_491_24;
  assign _GEN_136 = _T_532 ? _T_558 : _T_491_25;
  assign _GEN_137 = _T_532 ? _T_559 : _T_491_26;
  assign _GEN_138 = _T_532 ? _T_560 : _T_491_27;
  assign _GEN_139 = _T_532 ? _T_561 : _T_491_28;
  assign _GEN_140 = _T_532 ? _T_562 : _T_491_29;
  assign _GEN_141 = _T_532 ? _T_563 : _T_491_30;
  assign _GEN_142 = _T_532 ? _T_564 : _T_491_31;
  assign _GEN_143 = _T_532 ? 1'h1 : _T_531;
  assign _T_570 = _T_528 == 5'h1f;
  assign _T_574 = _T_528 + 5'h1;
  assign _T_575 = _T_574[4:0];
  assign _GEN_144 = _T_570 ? 1'h0 : _GEN_143;
  assign _GEN_145 = _T_570 ? 5'h0 : _T_575;
  assign _GEN_146 = _T_531 ? _GEN_144 : _GEN_143;
  assign _GEN_147 = _T_531 ? _GEN_145 : _T_528;
  assign _GEN_148 = _T_242 ? cores_1_inputMemAddr : cores_0_inputMemAddr;
  assign _GEN_149 = _T_242 ? cores_1_inputMemAddrValid : cores_0_inputMemAddrValid;
  assign _GEN_154 = _T_242 ? cores_1_inputMemBlockReady : cores_0_inputMemBlockReady;
  assign _GEN_162 = _T_242 ? cores_1_inputFinished : cores_0_inputFinished;
  assign _T_678 = _T_242 ? io_inputMemAddrReadys_1 : 1'h0;
  assign _GEN_164 = 5'h1 == _T_528 ? _T_491_1 : _T_491_0;
  assign _GEN_165 = 5'h2 == _T_528 ? _T_491_2 : _GEN_164;
  assign _GEN_166 = 5'h3 == _T_528 ? _T_491_3 : _GEN_165;
  assign _GEN_167 = 5'h4 == _T_528 ? _T_491_4 : _GEN_166;
  assign _GEN_168 = 5'h5 == _T_528 ? _T_491_5 : _GEN_167;
  assign _GEN_169 = 5'h6 == _T_528 ? _T_491_6 : _GEN_168;
  assign _GEN_170 = 5'h7 == _T_528 ? _T_491_7 : _GEN_169;
  assign _GEN_171 = 5'h8 == _T_528 ? _T_491_8 : _GEN_170;
  assign _GEN_172 = 5'h9 == _T_528 ? _T_491_9 : _GEN_171;
  assign _GEN_173 = 5'ha == _T_528 ? _T_491_10 : _GEN_172;
  assign _GEN_174 = 5'hb == _T_528 ? _T_491_11 : _GEN_173;
  assign _GEN_175 = 5'hc == _T_528 ? _T_491_12 : _GEN_174;
  assign _GEN_176 = 5'hd == _T_528 ? _T_491_13 : _GEN_175;
  assign _GEN_177 = 5'he == _T_528 ? _T_491_14 : _GEN_176;
  assign _GEN_178 = 5'hf == _T_528 ? _T_491_15 : _GEN_177;
  assign _GEN_179 = 5'h10 == _T_528 ? _T_491_16 : _GEN_178;
  assign _GEN_180 = 5'h11 == _T_528 ? _T_491_17 : _GEN_179;
  assign _GEN_181 = 5'h12 == _T_528 ? _T_491_18 : _GEN_180;
  assign _GEN_182 = 5'h13 == _T_528 ? _T_491_19 : _GEN_181;
  assign _GEN_183 = 5'h14 == _T_528 ? _T_491_20 : _GEN_182;
  assign _GEN_184 = 5'h15 == _T_528 ? _T_491_21 : _GEN_183;
  assign _GEN_185 = 5'h16 == _T_528 ? _T_491_22 : _GEN_184;
  assign _GEN_186 = 5'h17 == _T_528 ? _T_491_23 : _GEN_185;
  assign _GEN_187 = 5'h18 == _T_528 ? _T_491_24 : _GEN_186;
  assign _GEN_188 = 5'h19 == _T_528 ? _T_491_25 : _GEN_187;
  assign _GEN_189 = 5'h1a == _T_528 ? _T_491_26 : _GEN_188;
  assign _GEN_190 = 5'h1b == _T_528 ? _T_491_27 : _GEN_189;
  assign _GEN_191 = 5'h1c == _T_528 ? _T_491_28 : _GEN_190;
  assign _GEN_192 = 5'h1d == _T_528 ? _T_491_29 : _GEN_191;
  assign _GEN_193 = 5'h1e == _T_528 ? _T_491_30 : _GEN_192;
  assign _GEN_194 = 5'h1f == _T_528 ? _T_491_31 : _GEN_193;
  assign _T_683 = _T_242 ? _T_531 : 1'h0;
  assign _T_719 = _GEN_9_inputFinished | _T_570;
  assign _T_724 = _T_242 + 1'h1;
  assign _T_725 = _T_724[0:0];
  assign _T_726 = _T_242 ? 1'h1 : _T_725;
  assign _GEN_195 = _T_719 ? _T_726 : _T_242;
  assign _GEN_203 = _T_245 ? cores_1_outputMemAddr : cores_0_outputMemAddr;
  assign _GEN_204 = _T_245 ? cores_1_outputMemAddrValid : cores_0_outputMemAddrValid;
  assign _GEN_206 = _T_245 ? cores_1_outputMemBlock : cores_0_outputMemBlock;
  assign _GEN_207 = _T_245 ? cores_1_outputMemIdx : cores_0_outputMemIdx;
  assign _GEN_208 = _T_245 ? cores_1_outputMemBlockValid : cores_0_outputMemBlockValid;
  assign _GEN_211 = _T_245 ? cores_1_outputFinished : cores_0_outputFinished;
  assign _T_835 = _GEN_10_outputMemIdx == 5'h1f;
  assign _T_836 = _GEN_11_outputMemBlockValid & _T_835;
  assign _GEN_212 = _T_836 ? 1'h1 : _T_767;
  assign _T_839 = _T_767 == 1'h0;
  assign _GEN_213 = 5'h0 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_0;
  assign _GEN_214 = 5'h1 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_1;
  assign _GEN_215 = 5'h2 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_2;
  assign _GEN_216 = 5'h3 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_3;
  assign _GEN_217 = 5'h4 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_4;
  assign _GEN_218 = 5'h5 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_5;
  assign _GEN_219 = 5'h6 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_6;
  assign _GEN_220 = 5'h7 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_7;
  assign _GEN_221 = 5'h8 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_8;
  assign _GEN_222 = 5'h9 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_9;
  assign _GEN_223 = 5'ha == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_10;
  assign _GEN_224 = 5'hb == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_11;
  assign _GEN_225 = 5'hc == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_12;
  assign _GEN_226 = 5'hd == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_13;
  assign _GEN_227 = 5'he == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_14;
  assign _GEN_228 = 5'hf == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_15;
  assign _GEN_229 = 5'h10 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_16;
  assign _GEN_230 = 5'h11 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_17;
  assign _GEN_231 = 5'h12 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_18;
  assign _GEN_232 = 5'h13 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_19;
  assign _GEN_233 = 5'h14 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_20;
  assign _GEN_234 = 5'h15 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_21;
  assign _GEN_235 = 5'h16 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_22;
  assign _GEN_236 = 5'h17 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_23;
  assign _GEN_237 = 5'h18 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_24;
  assign _GEN_238 = 5'h19 == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_25;
  assign _GEN_239 = 5'h1a == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_26;
  assign _GEN_240 = 5'h1b == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_27;
  assign _GEN_241 = 5'h1c == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_28;
  assign _GEN_242 = 5'h1d == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_29;
  assign _GEN_243 = 5'h1e == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_30;
  assign _GEN_244 = 5'h1f == _GEN_12_outputMemIdx ? _GEN_13 : _T_730_31;
  assign _GEN_245 = _T_839 ? _GEN_213 : _T_730_0;
  assign _GEN_246 = _T_839 ? _GEN_214 : _T_730_1;
  assign _GEN_247 = _T_839 ? _GEN_215 : _T_730_2;
  assign _GEN_248 = _T_839 ? _GEN_216 : _T_730_3;
  assign _GEN_249 = _T_839 ? _GEN_217 : _T_730_4;
  assign _GEN_250 = _T_839 ? _GEN_218 : _T_730_5;
  assign _GEN_251 = _T_839 ? _GEN_219 : _T_730_6;
  assign _GEN_252 = _T_839 ? _GEN_220 : _T_730_7;
  assign _GEN_253 = _T_839 ? _GEN_221 : _T_730_8;
  assign _GEN_254 = _T_839 ? _GEN_222 : _T_730_9;
  assign _GEN_255 = _T_839 ? _GEN_223 : _T_730_10;
  assign _GEN_256 = _T_839 ? _GEN_224 : _T_730_11;
  assign _GEN_257 = _T_839 ? _GEN_225 : _T_730_12;
  assign _GEN_258 = _T_839 ? _GEN_226 : _T_730_13;
  assign _GEN_259 = _T_839 ? _GEN_227 : _T_730_14;
  assign _GEN_260 = _T_839 ? _GEN_228 : _T_730_15;
  assign _GEN_261 = _T_839 ? _GEN_229 : _T_730_16;
  assign _GEN_262 = _T_839 ? _GEN_230 : _T_730_17;
  assign _GEN_263 = _T_839 ? _GEN_231 : _T_730_18;
  assign _GEN_264 = _T_839 ? _GEN_232 : _T_730_19;
  assign _GEN_265 = _T_839 ? _GEN_233 : _T_730_20;
  assign _GEN_266 = _T_839 ? _GEN_234 : _T_730_21;
  assign _GEN_267 = _T_839 ? _GEN_235 : _T_730_22;
  assign _GEN_268 = _T_839 ? _GEN_236 : _T_730_23;
  assign _GEN_269 = _T_839 ? _GEN_237 : _T_730_24;
  assign _GEN_270 = _T_839 ? _GEN_238 : _T_730_25;
  assign _GEN_271 = _T_839 ? _GEN_239 : _T_730_26;
  assign _GEN_272 = _T_839 ? _GEN_240 : _T_730_27;
  assign _GEN_273 = _T_839 ? _GEN_241 : _T_730_28;
  assign _GEN_274 = _T_839 ? _GEN_242 : _T_730_29;
  assign _GEN_275 = _T_839 ? _GEN_243 : _T_730_30;
  assign _GEN_276 = _T_839 ? _GEN_244 : _T_730_31;
  assign _T_973 = {_T_730_1,_T_730_0};
  assign _T_974 = {_T_730_3,_T_730_2};
  assign _T_975 = {_T_974,_T_973};
  assign _T_976 = {_T_730_5,_T_730_4};
  assign _T_977 = {_T_730_7,_T_730_6};
  assign _T_978 = {_T_977,_T_976};
  assign _T_979 = {_T_978,_T_975};
  assign _T_980 = {_T_730_9,_T_730_8};
  assign _T_981 = {_T_730_11,_T_730_10};
  assign _T_982 = {_T_981,_T_980};
  assign _T_983 = {_T_730_13,_T_730_12};
  assign _T_984 = {_T_730_15,_T_730_14};
  assign _T_985 = {_T_984,_T_983};
  assign _T_986 = {_T_985,_T_982};
  assign _T_987 = {_T_986,_T_979};
  assign _T_988 = {_T_730_17,_T_730_16};
  assign _T_989 = {_T_730_19,_T_730_18};
  assign _T_990 = {_T_989,_T_988};
  assign _T_991 = {_T_730_21,_T_730_20};
  assign _T_992 = {_T_730_23,_T_730_22};
  assign _T_993 = {_T_992,_T_991};
  assign _T_994 = {_T_993,_T_990};
  assign _T_995 = {_T_730_25,_T_730_24};
  assign _T_996 = {_T_730_27,_T_730_26};
  assign _T_997 = {_T_996,_T_995};
  assign _T_998 = {_T_730_29,_T_730_28};
  assign _T_999 = {_T_730_31,_T_730_30};
  assign _T_1000 = {_T_999,_T_998};
  assign _T_1001 = {_T_1000,_T_997};
  assign _T_1002 = {_T_1001,_T_994};
  assign _T_1003 = {_T_1002,_T_987};
  assign _T_1005 = _T_245 == 1'h0;
  assign _T_1007 = _T_1005 ? io_outputMemAddrReadys_0 : 1'h0;
  assign _T_1010 = io_outputMemBlockReadys_0 & _T_767;
  assign _T_1012 = _T_1005 ? _T_1010 : 1'h0;
  assign _T_1013 = io_outputMemBlockReadys_0 & io_outputMemBlockValids_0;
  assign _T_1051 = _GEN_17_outputFinished | _T_1010;
  assign _T_1056 = _T_245 + 1'h1;
  assign _T_1057 = _T_1056[0:0];
  assign _T_1058 = _T_1005 ? 1'h0 : _T_1057;
  assign _GEN_277 = _T_1051 ? _T_1058 : _T_245;
  assign _GEN_278 = _T_1051 ? 1'h0 : _GEN_212;
  assign _GEN_286 = _T_248 ? cores_1_outputMemAddr : cores_0_outputMemAddr;
  assign _GEN_287 = _T_248 ? cores_1_outputMemAddrValid : cores_0_outputMemAddrValid;
  assign _GEN_289 = _T_248 ? cores_1_outputMemBlock : cores_0_outputMemBlock;
  assign _GEN_290 = _T_248 ? cores_1_outputMemIdx : cores_0_outputMemIdx;
  assign _GEN_291 = _T_248 ? cores_1_outputMemBlockValid : cores_0_outputMemBlockValid;
  assign _GEN_294 = _T_248 ? cores_1_outputFinished : cores_0_outputFinished;
  assign _T_1168 = _GEN_18_outputMemIdx == 5'h1f;
  assign _T_1169 = _GEN_19_outputMemBlockValid & _T_1168;
  assign _GEN_295 = _T_1169 ? 1'h1 : _T_1100;
  assign _T_1172 = _T_1100 == 1'h0;
  assign _GEN_296 = 5'h0 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_0;
  assign _GEN_297 = 5'h1 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_1;
  assign _GEN_298 = 5'h2 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_2;
  assign _GEN_299 = 5'h3 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_3;
  assign _GEN_300 = 5'h4 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_4;
  assign _GEN_301 = 5'h5 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_5;
  assign _GEN_302 = 5'h6 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_6;
  assign _GEN_303 = 5'h7 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_7;
  assign _GEN_304 = 5'h8 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_8;
  assign _GEN_305 = 5'h9 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_9;
  assign _GEN_306 = 5'ha == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_10;
  assign _GEN_307 = 5'hb == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_11;
  assign _GEN_308 = 5'hc == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_12;
  assign _GEN_309 = 5'hd == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_13;
  assign _GEN_310 = 5'he == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_14;
  assign _GEN_311 = 5'hf == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_15;
  assign _GEN_312 = 5'h10 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_16;
  assign _GEN_313 = 5'h11 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_17;
  assign _GEN_314 = 5'h12 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_18;
  assign _GEN_315 = 5'h13 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_19;
  assign _GEN_316 = 5'h14 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_20;
  assign _GEN_317 = 5'h15 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_21;
  assign _GEN_318 = 5'h16 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_22;
  assign _GEN_319 = 5'h17 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_23;
  assign _GEN_320 = 5'h18 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_24;
  assign _GEN_321 = 5'h19 == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_25;
  assign _GEN_322 = 5'h1a == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_26;
  assign _GEN_323 = 5'h1b == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_27;
  assign _GEN_324 = 5'h1c == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_28;
  assign _GEN_325 = 5'h1d == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_29;
  assign _GEN_326 = 5'h1e == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_30;
  assign _GEN_327 = 5'h1f == _GEN_20_outputMemIdx ? _GEN_21 : _T_1063_31;
  assign _GEN_328 = _T_1172 ? _GEN_296 : _T_1063_0;
  assign _GEN_329 = _T_1172 ? _GEN_297 : _T_1063_1;
  assign _GEN_330 = _T_1172 ? _GEN_298 : _T_1063_2;
  assign _GEN_331 = _T_1172 ? _GEN_299 : _T_1063_3;
  assign _GEN_332 = _T_1172 ? _GEN_300 : _T_1063_4;
  assign _GEN_333 = _T_1172 ? _GEN_301 : _T_1063_5;
  assign _GEN_334 = _T_1172 ? _GEN_302 : _T_1063_6;
  assign _GEN_335 = _T_1172 ? _GEN_303 : _T_1063_7;
  assign _GEN_336 = _T_1172 ? _GEN_304 : _T_1063_8;
  assign _GEN_337 = _T_1172 ? _GEN_305 : _T_1063_9;
  assign _GEN_338 = _T_1172 ? _GEN_306 : _T_1063_10;
  assign _GEN_339 = _T_1172 ? _GEN_307 : _T_1063_11;
  assign _GEN_340 = _T_1172 ? _GEN_308 : _T_1063_12;
  assign _GEN_341 = _T_1172 ? _GEN_309 : _T_1063_13;
  assign _GEN_342 = _T_1172 ? _GEN_310 : _T_1063_14;
  assign _GEN_343 = _T_1172 ? _GEN_311 : _T_1063_15;
  assign _GEN_344 = _T_1172 ? _GEN_312 : _T_1063_16;
  assign _GEN_345 = _T_1172 ? _GEN_313 : _T_1063_17;
  assign _GEN_346 = _T_1172 ? _GEN_314 : _T_1063_18;
  assign _GEN_347 = _T_1172 ? _GEN_315 : _T_1063_19;
  assign _GEN_348 = _T_1172 ? _GEN_316 : _T_1063_20;
  assign _GEN_349 = _T_1172 ? _GEN_317 : _T_1063_21;
  assign _GEN_350 = _T_1172 ? _GEN_318 : _T_1063_22;
  assign _GEN_351 = _T_1172 ? _GEN_319 : _T_1063_23;
  assign _GEN_352 = _T_1172 ? _GEN_320 : _T_1063_24;
  assign _GEN_353 = _T_1172 ? _GEN_321 : _T_1063_25;
  assign _GEN_354 = _T_1172 ? _GEN_322 : _T_1063_26;
  assign _GEN_355 = _T_1172 ? _GEN_323 : _T_1063_27;
  assign _GEN_356 = _T_1172 ? _GEN_324 : _T_1063_28;
  assign _GEN_357 = _T_1172 ? _GEN_325 : _T_1063_29;
  assign _GEN_358 = _T_1172 ? _GEN_326 : _T_1063_30;
  assign _GEN_359 = _T_1172 ? _GEN_327 : _T_1063_31;
  assign _T_1306 = {_T_1063_1,_T_1063_0};
  assign _T_1307 = {_T_1063_3,_T_1063_2};
  assign _T_1308 = {_T_1307,_T_1306};
  assign _T_1309 = {_T_1063_5,_T_1063_4};
  assign _T_1310 = {_T_1063_7,_T_1063_6};
  assign _T_1311 = {_T_1310,_T_1309};
  assign _T_1312 = {_T_1311,_T_1308};
  assign _T_1313 = {_T_1063_9,_T_1063_8};
  assign _T_1314 = {_T_1063_11,_T_1063_10};
  assign _T_1315 = {_T_1314,_T_1313};
  assign _T_1316 = {_T_1063_13,_T_1063_12};
  assign _T_1317 = {_T_1063_15,_T_1063_14};
  assign _T_1318 = {_T_1317,_T_1316};
  assign _T_1319 = {_T_1318,_T_1315};
  assign _T_1320 = {_T_1319,_T_1312};
  assign _T_1321 = {_T_1063_17,_T_1063_16};
  assign _T_1322 = {_T_1063_19,_T_1063_18};
  assign _T_1323 = {_T_1322,_T_1321};
  assign _T_1324 = {_T_1063_21,_T_1063_20};
  assign _T_1325 = {_T_1063_23,_T_1063_22};
  assign _T_1326 = {_T_1325,_T_1324};
  assign _T_1327 = {_T_1326,_T_1323};
  assign _T_1328 = {_T_1063_25,_T_1063_24};
  assign _T_1329 = {_T_1063_27,_T_1063_26};
  assign _T_1330 = {_T_1329,_T_1328};
  assign _T_1331 = {_T_1063_29,_T_1063_28};
  assign _T_1332 = {_T_1063_31,_T_1063_30};
  assign _T_1333 = {_T_1332,_T_1331};
  assign _T_1334 = {_T_1333,_T_1330};
  assign _T_1335 = {_T_1334,_T_1327};
  assign _T_1336 = {_T_1335,_T_1320};
  assign _T_1340 = _T_248 ? io_outputMemAddrReadys_1 : 1'h0;
  assign _T_1343 = io_outputMemBlockReadys_1 & _T_1100;
  assign _T_1345 = _T_248 ? _T_1343 : 1'h0;
  assign _T_1346 = io_outputMemBlockReadys_1 & io_outputMemBlockValids_1;
  assign _T_1384 = _GEN_25_outputFinished | _T_1343;
  assign _T_1389 = _T_248 + 1'h1;
  assign _T_1390 = _T_1389[0:0];
  assign _T_1391 = _T_248 ? 1'h1 : _T_1390;
  assign _GEN_360 = _T_1384 ? _T_1391 : _T_248;
  assign _GEN_361 = _T_1384 ? 1'h0 : _GEN_295;
  assign cumFinished = cores_0_outputFinished & cores_1_outputFinished;
  assign io_inputMemAddrs_0 = _GEN_0_inputMemAddr;
  assign io_inputMemAddrs_1 = _GEN_5_inputMemAddr;
  assign io_inputMemAddrValids_0 = _GEN_1_inputMemAddrValid;
  assign io_inputMemAddrValids_1 = _GEN_6_inputMemAddrValid;
  assign io_inputMemBlockReadys_0 = _GEN_2_inputMemBlockReady;
  assign io_inputMemBlockReadys_1 = _GEN_7_inputMemBlockReady;
  assign io_outputMemAddrs_0 = _GEN_15_outputMemAddr;
  assign io_outputMemAddrs_1 = _GEN_23_outputMemAddr;
  assign io_outputMemAddrValids_0 = _GEN_16_outputMemAddrValid;
  assign io_outputMemAddrValids_1 = _GEN_24_outputMemAddrValid;
  assign io_outputMemBlocks_0 = _T_1003;
  assign io_outputMemBlocks_1 = _T_1336;
  assign io_outputMemBlockValids_0 = _T_767;
  assign io_outputMemBlockValids_1 = _T_1100;
  assign io_finished = cumFinished;
  assign StreamingCore_io_inputMemAddrReady = cores_0_inputMemAddrReady;
  assign StreamingCore_io_inputMemBlock = cores_0_inputMemBlock;
  assign StreamingCore_io_inputMemIdx = cores_0_inputMemIdx;
  assign StreamingCore_io_inputMemBlockValid = cores_0_inputMemBlockValid;
  assign StreamingCore_io_outputMemAddrReady = cores_0_outputMemAddrReady;
  assign StreamingCore_io_outputMemBlockReady = cores_0_outputMemBlockReady;
  assign StreamingCore_clock = clock;
  assign StreamingCore_reset = reset;
  assign StreamingCore_1_io_inputMemAddrReady = cores_1_inputMemAddrReady;
  assign StreamingCore_1_io_inputMemBlock = cores_1_inputMemBlock;
  assign StreamingCore_1_io_inputMemIdx = cores_1_inputMemIdx;
  assign StreamingCore_1_io_inputMemBlockValid = cores_1_inputMemBlockValid;
  assign StreamingCore_1_io_outputMemAddrReady = cores_1_outputMemAddrReady;
  assign StreamingCore_1_io_outputMemBlockReady = cores_1_outputMemBlockReady;
  assign StreamingCore_1_clock = clock;
  assign StreamingCore_1_reset = reset;
  assign cores_0_inputMemAddr = StreamingCore_io_inputMemAddr;
  assign cores_0_inputMemAddrValid = StreamingCore_io_inputMemAddrValid;
  assign cores_0_inputMemAddrReady = _T_439;
  assign cores_0_inputMemBlock = _GEN_3;
  assign cores_0_inputMemIdx = _T_289;
  assign cores_0_inputMemBlockValid = _T_444;
  assign cores_0_inputMemBlockReady = StreamingCore_io_inputMemBlockReady;
  assign cores_0_outputMemAddr = StreamingCore_io_outputMemAddr;
  assign cores_0_outputMemAddrValid = StreamingCore_io_outputMemAddrValid;
  assign cores_0_outputMemAddrReady = _T_1007;
  assign cores_0_outputMemBlock = StreamingCore_io_outputMemBlock;
  assign cores_0_outputMemIdx = StreamingCore_io_outputMemIdx;
  assign cores_0_outputMemBlockValid = StreamingCore_io_outputMemBlockValid;
  assign cores_0_outputMemBlockReady = _T_1012;
  assign cores_0_inputFinished = StreamingCore_io_inputFinished;
  assign cores_0_outputFinished = StreamingCore_io_outputFinished;
  assign cores_1_inputMemAddr = StreamingCore_1_io_inputMemAddr;
  assign cores_1_inputMemAddrValid = StreamingCore_1_io_inputMemAddrValid;
  assign cores_1_inputMemAddrReady = _T_678;
  assign cores_1_inputMemBlock = _GEN_8;
  assign cores_1_inputMemIdx = _T_528;
  assign cores_1_inputMemBlockValid = _T_683;
  assign cores_1_inputMemBlockReady = StreamingCore_1_io_inputMemBlockReady;
  assign cores_1_outputMemAddr = StreamingCore_1_io_outputMemAddr;
  assign cores_1_outputMemAddrValid = StreamingCore_1_io_outputMemAddrValid;
  assign cores_1_outputMemAddrReady = _T_1340;
  assign cores_1_outputMemBlock = StreamingCore_1_io_outputMemBlock;
  assign cores_1_outputMemIdx = StreamingCore_1_io_outputMemIdx;
  assign cores_1_outputMemBlockValid = StreamingCore_1_io_outputMemBlockValid;
  assign cores_1_outputMemBlockReady = _T_1345;
  assign cores_1_inputFinished = StreamingCore_1_io_inputFinished;
  assign cores_1_outputFinished = StreamingCore_1_io_outputFinished;
  assign _GEN_0_inputMemAddr = _GEN_63;
  assign _GEN_1_inputMemAddrValid = _GEN_64;
  assign _GEN_2_inputMemBlockReady = _GEN_69;
  assign _GEN_3 = _GEN_109;
  assign _GEN_4_inputFinished = _GEN_77;
  assign _GEN_5_inputMemAddr = _GEN_148;
  assign _GEN_6_inputMemAddrValid = _GEN_149;
  assign _GEN_7_inputMemBlockReady = _GEN_154;
  assign _GEN_8 = _GEN_194;
  assign _GEN_9_inputFinished = _GEN_162;
  assign _GEN_10_outputMemIdx = _GEN_207;
  assign _GEN_11_outputMemBlockValid = _GEN_208;
  assign _GEN_12_outputMemIdx = _GEN_207;
  assign _GEN_13 = _GEN_14_outputMemBlock;
  assign _GEN_14_outputMemBlock = _GEN_206;
  assign _GEN_15_outputMemAddr = _GEN_203;
  assign _GEN_16_outputMemAddrValid = _GEN_204;
  assign _GEN_17_outputFinished = _GEN_211;
  assign _GEN_18_outputMemIdx = _GEN_290;
  assign _GEN_19_outputMemBlockValid = _GEN_291;
  assign _GEN_20_outputMemIdx = _GEN_290;
  assign _GEN_21 = _GEN_22_outputMemBlock;
  assign _GEN_22_outputMemBlock = _GEN_289;
  assign _GEN_23_outputMemAddr = _GEN_286;
  assign _GEN_24_outputMemAddrValid = _GEN_287;
  assign _GEN_25_outputFinished = _GEN_294;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_239 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_242 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_245 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_248 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_252_0 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_252_1 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_252_2 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_252_3 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_252_4 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_252_5 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_252_6 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_252_7 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_252_8 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_252_9 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_252_10 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_252_11 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_252_12 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_252_13 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_252_14 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_252_15 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_252_16 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_252_17 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_252_18 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_252_19 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_252_20 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_252_21 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_252_22 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_252_23 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_252_24 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_252_25 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_252_26 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_252_27 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_252_28 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_252_29 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_252_30 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_252_31 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_289 = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_292 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_491_0 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_491_1 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_491_2 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_491_3 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_491_4 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_491_5 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_491_6 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_491_7 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_491_8 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_491_9 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_491_10 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_491_11 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_491_12 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_491_13 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_491_14 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_491_15 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_491_16 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_491_17 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_491_18 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_491_19 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_491_20 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_491_21 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_491_22 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_491_23 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_491_24 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_491_25 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_491_26 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_491_27 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_491_28 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_491_29 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_491_30 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_491_31 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_528 = _RAND_70[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_531 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_730_0 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_730_1 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_730_2 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_730_3 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_730_4 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_730_5 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_730_6 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_730_7 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_730_8 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_730_9 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_730_10 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_730_11 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_730_12 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_730_13 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_730_14 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_730_15 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_730_16 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_730_17 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_730_18 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_730_19 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_730_20 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_730_21 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_730_22 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_730_23 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_730_24 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_730_25 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_730_26 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_730_27 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_730_28 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_730_29 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_730_30 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_730_31 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_767 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_1063_0 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_1063_1 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_1063_2 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_1063_3 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_1063_4 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_1063_5 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_1063_6 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_1063_7 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_1063_8 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_1063_9 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_1063_10 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_1063_11 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_1063_12 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_1063_13 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_1063_14 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_1063_15 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_1063_16 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_1063_17 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_1063_18 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_1063_19 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_1063_20 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_1063_21 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_1063_22 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_1063_23 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_1063_24 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_1063_25 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_1063_26 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_1063_27 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_1063_28 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_1063_29 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  _T_1063_30 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_1063_31 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  _T_1100 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      if (_T_480) begin
        if (_T_437) begin
          _T_239 <= 1'h0;
        end else begin
          _T_239 <= _T_486;
        end
      end
    end
    if (reset) begin
      _T_242 <= 1'h1;
    end else begin
      if (_T_719) begin
        if (_T_242) begin
          _T_242 <= 1'h1;
        end else begin
          _T_242 <= _T_725;
        end
      end
    end
    if (reset) begin
      _T_245 <= 1'h0;
    end else begin
      if (_T_1051) begin
        if (_T_1005) begin
          _T_245 <= 1'h0;
        end else begin
          _T_245 <= _T_1057;
        end
      end
    end
    if (reset) begin
      _T_248 <= 1'h1;
    end else begin
      if (_T_1384) begin
        if (_T_248) begin
          _T_248 <= 1'h1;
        end else begin
          _T_248 <= _T_1390;
        end
      end
    end
    if (_T_293) begin
      _T_252_0 <= _T_294;
    end
    if (_T_293) begin
      _T_252_1 <= _T_295;
    end
    if (_T_293) begin
      _T_252_2 <= _T_296;
    end
    if (_T_293) begin
      _T_252_3 <= _T_297;
    end
    if (_T_293) begin
      _T_252_4 <= _T_298;
    end
    if (_T_293) begin
      _T_252_5 <= _T_299;
    end
    if (_T_293) begin
      _T_252_6 <= _T_300;
    end
    if (_T_293) begin
      _T_252_7 <= _T_301;
    end
    if (_T_293) begin
      _T_252_8 <= _T_302;
    end
    if (_T_293) begin
      _T_252_9 <= _T_303;
    end
    if (_T_293) begin
      _T_252_10 <= _T_304;
    end
    if (_T_293) begin
      _T_252_11 <= _T_305;
    end
    if (_T_293) begin
      _T_252_12 <= _T_306;
    end
    if (_T_293) begin
      _T_252_13 <= _T_307;
    end
    if (_T_293) begin
      _T_252_14 <= _T_308;
    end
    if (_T_293) begin
      _T_252_15 <= _T_309;
    end
    if (_T_293) begin
      _T_252_16 <= _T_310;
    end
    if (_T_293) begin
      _T_252_17 <= _T_311;
    end
    if (_T_293) begin
      _T_252_18 <= _T_312;
    end
    if (_T_293) begin
      _T_252_19 <= _T_313;
    end
    if (_T_293) begin
      _T_252_20 <= _T_314;
    end
    if (_T_293) begin
      _T_252_21 <= _T_315;
    end
    if (_T_293) begin
      _T_252_22 <= _T_316;
    end
    if (_T_293) begin
      _T_252_23 <= _T_317;
    end
    if (_T_293) begin
      _T_252_24 <= _T_318;
    end
    if (_T_293) begin
      _T_252_25 <= _T_319;
    end
    if (_T_293) begin
      _T_252_26 <= _T_320;
    end
    if (_T_293) begin
      _T_252_27 <= _T_321;
    end
    if (_T_293) begin
      _T_252_28 <= _T_322;
    end
    if (_T_293) begin
      _T_252_29 <= _T_323;
    end
    if (_T_293) begin
      _T_252_30 <= _T_324;
    end
    if (_T_293) begin
      _T_252_31 <= _T_325;
    end
    if (reset) begin
      _T_289 <= 5'h0;
    end else begin
      if (_T_292) begin
        if (_T_331) begin
          _T_289 <= 5'h0;
        end else begin
          _T_289 <= _T_336;
        end
      end
    end
    if (reset) begin
      _T_292 <= 1'h0;
    end else begin
      if (_T_292) begin
        if (_T_331) begin
          _T_292 <= 1'h0;
        end else begin
          if (_T_293) begin
            _T_292 <= 1'h1;
          end
        end
      end else begin
        if (_T_293) begin
          _T_292 <= 1'h1;
        end
      end
    end
    if (_T_532) begin
      _T_491_0 <= _T_533;
    end
    if (_T_532) begin
      _T_491_1 <= _T_534;
    end
    if (_T_532) begin
      _T_491_2 <= _T_535;
    end
    if (_T_532) begin
      _T_491_3 <= _T_536;
    end
    if (_T_532) begin
      _T_491_4 <= _T_537;
    end
    if (_T_532) begin
      _T_491_5 <= _T_538;
    end
    if (_T_532) begin
      _T_491_6 <= _T_539;
    end
    if (_T_532) begin
      _T_491_7 <= _T_540;
    end
    if (_T_532) begin
      _T_491_8 <= _T_541;
    end
    if (_T_532) begin
      _T_491_9 <= _T_542;
    end
    if (_T_532) begin
      _T_491_10 <= _T_543;
    end
    if (_T_532) begin
      _T_491_11 <= _T_544;
    end
    if (_T_532) begin
      _T_491_12 <= _T_545;
    end
    if (_T_532) begin
      _T_491_13 <= _T_546;
    end
    if (_T_532) begin
      _T_491_14 <= _T_547;
    end
    if (_T_532) begin
      _T_491_15 <= _T_548;
    end
    if (_T_532) begin
      _T_491_16 <= _T_549;
    end
    if (_T_532) begin
      _T_491_17 <= _T_550;
    end
    if (_T_532) begin
      _T_491_18 <= _T_551;
    end
    if (_T_532) begin
      _T_491_19 <= _T_552;
    end
    if (_T_532) begin
      _T_491_20 <= _T_553;
    end
    if (_T_532) begin
      _T_491_21 <= _T_554;
    end
    if (_T_532) begin
      _T_491_22 <= _T_555;
    end
    if (_T_532) begin
      _T_491_23 <= _T_556;
    end
    if (_T_532) begin
      _T_491_24 <= _T_557;
    end
    if (_T_532) begin
      _T_491_25 <= _T_558;
    end
    if (_T_532) begin
      _T_491_26 <= _T_559;
    end
    if (_T_532) begin
      _T_491_27 <= _T_560;
    end
    if (_T_532) begin
      _T_491_28 <= _T_561;
    end
    if (_T_532) begin
      _T_491_29 <= _T_562;
    end
    if (_T_532) begin
      _T_491_30 <= _T_563;
    end
    if (_T_532) begin
      _T_491_31 <= _T_564;
    end
    if (reset) begin
      _T_528 <= 5'h0;
    end else begin
      if (_T_531) begin
        if (_T_570) begin
          _T_528 <= 5'h0;
        end else begin
          _T_528 <= _T_575;
        end
      end
    end
    if (reset) begin
      _T_531 <= 1'h0;
    end else begin
      if (_T_531) begin
        if (_T_570) begin
          _T_531 <= 1'h0;
        end else begin
          if (_T_532) begin
            _T_531 <= 1'h1;
          end
        end
      end else begin
        if (_T_532) begin
          _T_531 <= 1'h1;
        end
      end
    end
    if (_T_839) begin
      if (5'h0 == _GEN_12_outputMemIdx) begin
        _T_730_0 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h1 == _GEN_12_outputMemIdx) begin
        _T_730_1 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h2 == _GEN_12_outputMemIdx) begin
        _T_730_2 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h3 == _GEN_12_outputMemIdx) begin
        _T_730_3 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h4 == _GEN_12_outputMemIdx) begin
        _T_730_4 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h5 == _GEN_12_outputMemIdx) begin
        _T_730_5 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h6 == _GEN_12_outputMemIdx) begin
        _T_730_6 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h7 == _GEN_12_outputMemIdx) begin
        _T_730_7 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h8 == _GEN_12_outputMemIdx) begin
        _T_730_8 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h9 == _GEN_12_outputMemIdx) begin
        _T_730_9 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'ha == _GEN_12_outputMemIdx) begin
        _T_730_10 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'hb == _GEN_12_outputMemIdx) begin
        _T_730_11 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'hc == _GEN_12_outputMemIdx) begin
        _T_730_12 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'hd == _GEN_12_outputMemIdx) begin
        _T_730_13 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'he == _GEN_12_outputMemIdx) begin
        _T_730_14 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'hf == _GEN_12_outputMemIdx) begin
        _T_730_15 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h10 == _GEN_12_outputMemIdx) begin
        _T_730_16 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h11 == _GEN_12_outputMemIdx) begin
        _T_730_17 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h12 == _GEN_12_outputMemIdx) begin
        _T_730_18 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h13 == _GEN_12_outputMemIdx) begin
        _T_730_19 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h14 == _GEN_12_outputMemIdx) begin
        _T_730_20 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h15 == _GEN_12_outputMemIdx) begin
        _T_730_21 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h16 == _GEN_12_outputMemIdx) begin
        _T_730_22 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h17 == _GEN_12_outputMemIdx) begin
        _T_730_23 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h18 == _GEN_12_outputMemIdx) begin
        _T_730_24 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h19 == _GEN_12_outputMemIdx) begin
        _T_730_25 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h1a == _GEN_12_outputMemIdx) begin
        _T_730_26 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h1b == _GEN_12_outputMemIdx) begin
        _T_730_27 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h1c == _GEN_12_outputMemIdx) begin
        _T_730_28 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h1d == _GEN_12_outputMemIdx) begin
        _T_730_29 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h1e == _GEN_12_outputMemIdx) begin
        _T_730_30 <= _GEN_13;
      end
    end
    if (_T_839) begin
      if (5'h1f == _GEN_12_outputMemIdx) begin
        _T_730_31 <= _GEN_13;
      end
    end
    if (reset) begin
      _T_767 <= 1'h0;
    end else begin
      if (_T_1051) begin
        _T_767 <= 1'h0;
      end else begin
        if (_T_836) begin
          _T_767 <= 1'h1;
        end
      end
    end
    if (_T_1172) begin
      if (5'h0 == _GEN_20_outputMemIdx) begin
        _T_1063_0 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h1 == _GEN_20_outputMemIdx) begin
        _T_1063_1 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h2 == _GEN_20_outputMemIdx) begin
        _T_1063_2 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h3 == _GEN_20_outputMemIdx) begin
        _T_1063_3 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h4 == _GEN_20_outputMemIdx) begin
        _T_1063_4 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h5 == _GEN_20_outputMemIdx) begin
        _T_1063_5 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h6 == _GEN_20_outputMemIdx) begin
        _T_1063_6 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h7 == _GEN_20_outputMemIdx) begin
        _T_1063_7 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h8 == _GEN_20_outputMemIdx) begin
        _T_1063_8 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h9 == _GEN_20_outputMemIdx) begin
        _T_1063_9 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'ha == _GEN_20_outputMemIdx) begin
        _T_1063_10 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'hb == _GEN_20_outputMemIdx) begin
        _T_1063_11 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'hc == _GEN_20_outputMemIdx) begin
        _T_1063_12 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'hd == _GEN_20_outputMemIdx) begin
        _T_1063_13 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'he == _GEN_20_outputMemIdx) begin
        _T_1063_14 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'hf == _GEN_20_outputMemIdx) begin
        _T_1063_15 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h10 == _GEN_20_outputMemIdx) begin
        _T_1063_16 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h11 == _GEN_20_outputMemIdx) begin
        _T_1063_17 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h12 == _GEN_20_outputMemIdx) begin
        _T_1063_18 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h13 == _GEN_20_outputMemIdx) begin
        _T_1063_19 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h14 == _GEN_20_outputMemIdx) begin
        _T_1063_20 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h15 == _GEN_20_outputMemIdx) begin
        _T_1063_21 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h16 == _GEN_20_outputMemIdx) begin
        _T_1063_22 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h17 == _GEN_20_outputMemIdx) begin
        _T_1063_23 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h18 == _GEN_20_outputMemIdx) begin
        _T_1063_24 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h19 == _GEN_20_outputMemIdx) begin
        _T_1063_25 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h1a == _GEN_20_outputMemIdx) begin
        _T_1063_26 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h1b == _GEN_20_outputMemIdx) begin
        _T_1063_27 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h1c == _GEN_20_outputMemIdx) begin
        _T_1063_28 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h1d == _GEN_20_outputMemIdx) begin
        _T_1063_29 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h1e == _GEN_20_outputMemIdx) begin
        _T_1063_30 <= _GEN_21;
      end
    end
    if (_T_1172) begin
      if (5'h1f == _GEN_20_outputMemIdx) begin
        _T_1063_31 <= _GEN_21;
      end
    end
    if (reset) begin
      _T_1100 <= 1'h0;
    end else begin
      if (_T_1384) begin
        _T_1100 <= 1'h0;
      end else begin
        if (_T_1169) begin
          _T_1100 <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_293 & _T_329) begin
          $fwrite(32'h80000002,"inputBuffer: 0x%h for core %d, channel 0\n",io_inputMemBlocks_0,_T_239);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_532 & _T_329) begin
          $fwrite(32'h80000002,"inputBuffer: 0x%h for core %d, channel 1\n",io_inputMemBlocks_1,_T_242);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1013 & _T_329) begin
          $fwrite(32'h80000002,"outputBuffer: 0x%h for core %d, channel 0\n",io_outputMemBlocks_0,_T_245);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1346 & _T_329) begin
          $fwrite(32'h80000002,"outputBuffer: 0x%h for core %d, channel 1\n",io_outputMemBlocks_1,_T_248);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
