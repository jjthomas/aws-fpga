`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module DualPortBRAM(
  input         clock,
  input  [4:0]  io_a_addr,
  input  [15:0] io_a_din,
  input         io_a_wr,
  input  [4:0]  io_b_addr,
  output [15:0] io_b_dout
);
  reg [15:0] mem [0:31];
  reg [31:0] _RAND_0;
  wire [15:0] mem__T_12_data;
  wire [4:0] mem__T_12_addr;
  wire [15:0] mem__T_14_data;
  wire [4:0] mem__T_14_addr;
  wire [15:0] mem__T_13_data;
  wire [4:0] mem__T_13_addr;
  wire  mem__T_13_mask;
  wire  mem__T_13_en;
  wire [15:0] mem__T_15_data;
  wire [4:0] mem__T_15_addr;
  wire  mem__T_15_mask;
  wire  mem__T_15_en;
  wire  _GEN_8;
  reg [4:0] mem__T_12_addr_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] mem__T_14_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign mem__T_12_addr = mem__T_12_addr_pipe_0;
  assign mem__T_12_data = mem[mem__T_12_addr];
  assign mem__T_14_addr = mem__T_14_addr_pipe_0;
  assign mem__T_14_data = mem[mem__T_14_addr];
  assign mem__T_13_data = io_a_din;
  assign mem__T_13_addr = io_a_addr;
  assign mem__T_13_mask = io_a_wr;
  assign mem__T_13_en = io_a_wr;
  assign mem__T_15_data = 16'h0;
  assign mem__T_15_addr = io_b_addr;
  assign mem__T_15_mask = 1'h0;
  assign mem__T_15_en = 1'h0;
  assign _GEN_8 = 1'h1;
  assign io_b_dout = mem__T_14_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem__T_12_addr_pipe_0 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem__T_14_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_13_en & mem__T_13_mask) begin
      mem[mem__T_13_addr] <= mem__T_13_data;
    end
    if(mem__T_15_en & mem__T_15_mask) begin
      mem[mem__T_15_addr] <= mem__T_15_data;
    end
    if (_GEN_8) begin
      mem__T_12_addr_pipe_0 <= io_a_addr;
    end
    if (_GEN_8) begin
      mem__T_14_addr_pipe_0 <= io_b_addr;
    end
  end
endmodule
module PassThrough(
  input         clock,
  input         reset,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  input  [9:0]  io_inputBits,
  output        io_inputMemConsumed,
  input         io_inputFinished,
  output [15:0] io_outputMemBlock,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output [9:0]  io_outputBits,
  output        io_outputFinished,
  input         io_outputMemFlushed
);
  reg  inputMemBlock_0;
  reg [31:0] _RAND_0;
  reg  inputMemBlock_1;
  reg [31:0] _RAND_1;
  reg  inputMemBlock_2;
  reg [31:0] _RAND_2;
  reg  inputMemBlock_3;
  reg [31:0] _RAND_3;
  reg  inputMemBlock_4;
  reg [31:0] _RAND_4;
  reg  inputMemBlock_5;
  reg [31:0] _RAND_5;
  reg  inputMemBlock_6;
  reg [31:0] _RAND_6;
  reg  inputMemBlock_7;
  reg [31:0] _RAND_7;
  reg  inputMemBlock_8;
  reg [31:0] _RAND_8;
  reg  inputMemBlock_9;
  reg [31:0] _RAND_9;
  reg  inputMemBlock_10;
  reg [31:0] _RAND_10;
  reg  inputMemBlock_11;
  reg [31:0] _RAND_11;
  reg  inputMemBlock_12;
  reg [31:0] _RAND_12;
  reg  inputMemBlock_13;
  reg [31:0] _RAND_13;
  reg  inputMemBlock_14;
  reg [31:0] _RAND_14;
  reg  inputMemBlock_15;
  reg [31:0] _RAND_15;
  reg [4:0] inputPieceBitsRemaining;
  reg [31:0] _RAND_16;
  reg [9:0] inputBitsRemaining;
  reg [31:0] _RAND_17;
  reg  inputBlockLoaded;
  reg [31:0] _RAND_18;
  reg  outputMemBlock_0;
  reg [31:0] _RAND_19;
  reg  outputMemBlock_1;
  reg [31:0] _RAND_20;
  reg  outputMemBlock_2;
  reg [31:0] _RAND_21;
  reg  outputMemBlock_3;
  reg [31:0] _RAND_22;
  reg  outputMemBlock_4;
  reg [31:0] _RAND_23;
  reg  outputMemBlock_5;
  reg [31:0] _RAND_24;
  reg  outputMemBlock_6;
  reg [31:0] _RAND_25;
  reg  outputMemBlock_7;
  reg [31:0] _RAND_26;
  reg  outputMemBlock_8;
  reg [31:0] _RAND_27;
  reg  outputMemBlock_9;
  reg [31:0] _RAND_28;
  reg  outputMemBlock_10;
  reg [31:0] _RAND_29;
  reg  outputMemBlock_11;
  reg [31:0] _RAND_30;
  reg  outputMemBlock_12;
  reg [31:0] _RAND_31;
  reg  outputMemBlock_13;
  reg [31:0] _RAND_32;
  reg  outputMemBlock_14;
  reg [31:0] _RAND_33;
  reg  outputMemBlock_15;
  reg [31:0] _RAND_34;
  reg [9:0] outputBits;
  reg [31:0] _RAND_35;
  reg [4:0] outputPieceBits;
  reg [31:0] _RAND_36;
  wire  inputBram_clock;
  wire [4:0] inputBram_io_a_addr;
  wire [15:0] inputBram_io_a_din;
  wire  inputBram_io_a_wr;
  wire [4:0] inputBram_io_b_addr;
  wire [15:0] inputBram_io_b_dout;
  reg [4:0] inputReadAddr;
  reg [31:0] _RAND_37;
  reg  inputPieceRead;
  reg [31:0] _RAND_38;
  wire  outputBram_clock;
  wire [4:0] outputBram_io_a_addr;
  wire [15:0] outputBram_io_a_din;
  wire  outputBram_io_a_wr;
  wire [4:0] outputBram_io_b_addr;
  wire [15:0] outputBram_io_b_dout;
  reg [4:0] outputWriteAddr;
  reg [31:0] _RAND_39;
  reg [4:0] outputReadAddr;
  reg [31:0] _RAND_40;
  wire  _T_75;
  wire  _T_76;
  wire  _GEN_0;
  wire [9:0] _GEN_1;
  wire  _T_79;
  wire  _T_80;
  wire  _GEN_2;
  wire  _T_84;
  wire  _T_85;
  wire  _T_89;
  wire  _T_90;
  wire  _T_92;
  wire  _T_96;
  wire [9:0] _T_98;
  wire [5:0] _T_100;
  wire [4:0] _T_101;
  wire  _T_102;
  wire  _T_103;
  wire  _T_104;
  wire  _T_105;
  wire  _T_106;
  wire  _T_107;
  wire  _T_108;
  wire  _T_109;
  wire  _T_110;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  _T_114;
  wire  _T_115;
  wire  _T_116;
  wire  _T_117;
  wire [9:0] _GEN_4;
  wire [4:0] _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [9:0] _GEN_23;
  wire [4:0] _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  inputAdvance;
  wire  _T_120;
  wire  _T_122;
  wire  _T_124;
  wire  _T_125;
  wire  _T_129;
  wire  _T_130;
  wire [5:0] _T_132;
  wire [5:0] _T_133;
  wire [4:0] _T_134;
  wire [10:0] _T_136;
  wire [10:0] _T_137;
  wire [9:0] _T_138;
  wire [9:0] _GEN_41;
  wire [9:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  nextBitValid;
  wire  nextBit;
  wire [5:0] _T_142;
  wire [4:0] _T_143;
  wire [10:0] _T_145;
  wire [9:0] _T_146;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire [4:0] _GEN_74;
  wire [9:0] _GEN_75;
  wire  _T_148;
  wire  _T_151;
  wire  _T_153;
  wire  _T_154;
  wire  _T_155;
  wire [1:0] _T_156;
  wire [1:0] _T_157;
  wire [3:0] _T_158;
  wire [1:0] _T_159;
  wire [1:0] _T_160;
  wire [3:0] _T_161;
  wire [7:0] _T_162;
  wire [1:0] _T_163;
  wire [1:0] _T_164;
  wire [3:0] _T_165;
  wire [1:0] _T_166;
  wire [1:0] _T_167;
  wire [3:0] _T_168;
  wire [7:0] _T_169;
  wire [15:0] _T_170;
  wire [5:0] _T_175;
  wire [4:0] _T_176;
  wire [4:0] _GEN_76;
  wire [4:0] _GEN_77;
  reg  outputReadingStarted;
  reg [31:0] _RAND_41;
  wire  _T_181;
  wire  _T_188;
  wire  _T_189;
  wire  _T_190;
  wire  _T_191;
  wire  _GEN_78;
  wire  _T_193;
  wire  _T_195;
  wire  _T_196;
  wire [5:0] _T_198;
  wire [4:0] _T_199;
  wire [4:0] _GEN_79;
  wire  _T_203;
  wire  _T_204;
  wire  _T_214;
  wire  _T_219;
  wire  _T_220;
  wire [9:0] _GEN_80;
  wire [4:0] _GEN_81;
  wire  _GEN_82;
  wire [4:0] _GEN_83;
  wire [4:0] _GEN_84;
  DualPortBRAM inputBram (
    .clock(inputBram_clock),
    .io_a_addr(inputBram_io_a_addr),
    .io_a_din(inputBram_io_a_din),
    .io_a_wr(inputBram_io_a_wr),
    .io_b_addr(inputBram_io_b_addr),
    .io_b_dout(inputBram_io_b_dout)
  );
  DualPortBRAM outputBram (
    .clock(outputBram_clock),
    .io_a_addr(outputBram_io_a_addr),
    .io_a_din(outputBram_io_a_din),
    .io_a_wr(outputBram_io_a_wr),
    .io_b_addr(outputBram_io_b_addr),
    .io_b_dout(outputBram_io_b_dout)
  );
  assign _T_75 = io_inputMemIdx == 5'h1f;
  assign _T_76 = io_inputMemBlockValid & _T_75;
  assign _GEN_0 = _T_76 ? 1'h1 : inputBlockLoaded;
  assign _GEN_1 = _T_76 ? io_inputBits : inputBitsRemaining;
  assign _T_79 = inputBitsRemaining == 10'h0;
  assign _T_80 = inputBlockLoaded & _T_79;
  assign _GEN_2 = _T_80 ? 1'h0 : _GEN_0;
  assign _T_84 = inputPieceBitsRemaining == 5'h0;
  assign _T_85 = inputBlockLoaded & _T_84;
  assign _T_89 = _T_79 == 1'h0;
  assign _T_90 = _T_85 & _T_89;
  assign _T_92 = inputPieceRead == 1'h0;
  assign _T_96 = inputBitsRemaining < 10'h10;
  assign _T_98 = _T_96 ? inputBitsRemaining : 10'h10;
  assign _T_100 = inputReadAddr + 5'h1;
  assign _T_101 = _T_100[4:0];
  assign _T_102 = inputBram_io_b_dout[0];
  assign _T_103 = inputBram_io_b_dout[1];
  assign _T_104 = inputBram_io_b_dout[2];
  assign _T_105 = inputBram_io_b_dout[3];
  assign _T_106 = inputBram_io_b_dout[4];
  assign _T_107 = inputBram_io_b_dout[5];
  assign _T_108 = inputBram_io_b_dout[6];
  assign _T_109 = inputBram_io_b_dout[7];
  assign _T_110 = inputBram_io_b_dout[8];
  assign _T_111 = inputBram_io_b_dout[9];
  assign _T_112 = inputBram_io_b_dout[10];
  assign _T_113 = inputBram_io_b_dout[11];
  assign _T_114 = inputBram_io_b_dout[12];
  assign _T_115 = inputBram_io_b_dout[13];
  assign _T_116 = inputBram_io_b_dout[14];
  assign _T_117 = inputBram_io_b_dout[15];
  assign _GEN_4 = _T_92 ? {{5'd0}, inputPieceBitsRemaining} : _T_98;
  assign _GEN_5 = _T_92 ? inputReadAddr : _T_101;
  assign _GEN_6 = _T_92 ? inputMemBlock_0 : _T_102;
  assign _GEN_7 = _T_92 ? inputMemBlock_1 : _T_103;
  assign _GEN_8 = _T_92 ? inputMemBlock_2 : _T_104;
  assign _GEN_9 = _T_92 ? inputMemBlock_3 : _T_105;
  assign _GEN_10 = _T_92 ? inputMemBlock_4 : _T_106;
  assign _GEN_11 = _T_92 ? inputMemBlock_5 : _T_107;
  assign _GEN_12 = _T_92 ? inputMemBlock_6 : _T_108;
  assign _GEN_13 = _T_92 ? inputMemBlock_7 : _T_109;
  assign _GEN_14 = _T_92 ? inputMemBlock_8 : _T_110;
  assign _GEN_15 = _T_92 ? inputMemBlock_9 : _T_111;
  assign _GEN_16 = _T_92 ? inputMemBlock_10 : _T_112;
  assign _GEN_17 = _T_92 ? inputMemBlock_11 : _T_113;
  assign _GEN_18 = _T_92 ? inputMemBlock_12 : _T_114;
  assign _GEN_19 = _T_92 ? inputMemBlock_13 : _T_115;
  assign _GEN_20 = _T_92 ? inputMemBlock_14 : _T_116;
  assign _GEN_21 = _T_92 ? inputMemBlock_15 : _T_117;
  assign _GEN_22 = _T_90 ? _T_92 : inputPieceRead;
  assign _GEN_23 = _T_90 ? _GEN_4 : {{5'd0}, inputPieceBitsRemaining};
  assign _GEN_24 = _T_90 ? _GEN_5 : inputReadAddr;
  assign _GEN_25 = _T_90 ? _GEN_6 : inputMemBlock_0;
  assign _GEN_26 = _T_90 ? _GEN_7 : inputMemBlock_1;
  assign _GEN_27 = _T_90 ? _GEN_8 : inputMemBlock_2;
  assign _GEN_28 = _T_90 ? _GEN_9 : inputMemBlock_3;
  assign _GEN_29 = _T_90 ? _GEN_10 : inputMemBlock_4;
  assign _GEN_30 = _T_90 ? _GEN_11 : inputMemBlock_5;
  assign _GEN_31 = _T_90 ? _GEN_12 : inputMemBlock_6;
  assign _GEN_32 = _T_90 ? _GEN_13 : inputMemBlock_7;
  assign _GEN_33 = _T_90 ? _GEN_14 : inputMemBlock_8;
  assign _GEN_34 = _T_90 ? _GEN_15 : inputMemBlock_9;
  assign _GEN_35 = _T_90 ? _GEN_16 : inputMemBlock_10;
  assign _GEN_36 = _T_90 ? _GEN_17 : inputMemBlock_11;
  assign _GEN_37 = _T_90 ? _GEN_18 : inputMemBlock_12;
  assign _GEN_38 = _T_90 ? _GEN_19 : inputMemBlock_13;
  assign _GEN_39 = _T_90 ? _GEN_20 : inputMemBlock_14;
  assign _GEN_40 = _T_90 ? _GEN_21 : inputMemBlock_15;
  assign _T_120 = outputPieceBits != 5'h10;
  assign _T_122 = outputBits == 10'h200;
  assign _T_124 = _T_122 == 1'h0;
  assign _T_125 = _T_120 & _T_124;
  assign _T_129 = _T_84 == 1'h0;
  assign _T_130 = _T_125 & _T_129;
  assign _T_132 = inputPieceBitsRemaining - 5'h1;
  assign _T_133 = $unsigned(_T_132);
  assign _T_134 = _T_133[4:0];
  assign _T_136 = inputBitsRemaining - 10'h1;
  assign _T_137 = $unsigned(_T_136);
  assign _T_138 = _T_137[9:0];
  assign _GEN_41 = inputAdvance ? {{5'd0}, _T_134} : _GEN_23;
  assign _GEN_42 = inputAdvance ? _T_138 : _GEN_1;
  assign _GEN_43 = inputAdvance ? inputMemBlock_1 : _GEN_25;
  assign _GEN_44 = inputAdvance ? inputMemBlock_2 : _GEN_26;
  assign _GEN_45 = inputAdvance ? inputMemBlock_3 : _GEN_27;
  assign _GEN_46 = inputAdvance ? inputMemBlock_4 : _GEN_28;
  assign _GEN_47 = inputAdvance ? inputMemBlock_5 : _GEN_29;
  assign _GEN_48 = inputAdvance ? inputMemBlock_6 : _GEN_30;
  assign _GEN_49 = inputAdvance ? inputMemBlock_7 : _GEN_31;
  assign _GEN_50 = inputAdvance ? inputMemBlock_8 : _GEN_32;
  assign _GEN_51 = inputAdvance ? inputMemBlock_9 : _GEN_33;
  assign _GEN_52 = inputAdvance ? inputMemBlock_10 : _GEN_34;
  assign _GEN_53 = inputAdvance ? inputMemBlock_11 : _GEN_35;
  assign _GEN_54 = inputAdvance ? inputMemBlock_12 : _GEN_36;
  assign _GEN_55 = inputAdvance ? inputMemBlock_13 : _GEN_37;
  assign _GEN_56 = inputAdvance ? inputMemBlock_14 : _GEN_38;
  assign _GEN_57 = inputAdvance ? inputMemBlock_15 : _GEN_39;
  assign _T_142 = outputPieceBits + 5'h1;
  assign _T_143 = _T_142[4:0];
  assign _T_145 = outputBits + 10'h1;
  assign _T_146 = _T_145[9:0];
  assign _GEN_58 = nextBitValid ? nextBit : outputMemBlock_15;
  assign _GEN_59 = nextBitValid ? outputMemBlock_1 : outputMemBlock_0;
  assign _GEN_60 = nextBitValid ? outputMemBlock_2 : outputMemBlock_1;
  assign _GEN_61 = nextBitValid ? outputMemBlock_3 : outputMemBlock_2;
  assign _GEN_62 = nextBitValid ? outputMemBlock_4 : outputMemBlock_3;
  assign _GEN_63 = nextBitValid ? outputMemBlock_5 : outputMemBlock_4;
  assign _GEN_64 = nextBitValid ? outputMemBlock_6 : outputMemBlock_5;
  assign _GEN_65 = nextBitValid ? outputMemBlock_7 : outputMemBlock_6;
  assign _GEN_66 = nextBitValid ? outputMemBlock_8 : outputMemBlock_7;
  assign _GEN_67 = nextBitValid ? outputMemBlock_9 : outputMemBlock_8;
  assign _GEN_68 = nextBitValid ? outputMemBlock_10 : outputMemBlock_9;
  assign _GEN_69 = nextBitValid ? outputMemBlock_11 : outputMemBlock_10;
  assign _GEN_70 = nextBitValid ? outputMemBlock_12 : outputMemBlock_11;
  assign _GEN_71 = nextBitValid ? outputMemBlock_13 : outputMemBlock_12;
  assign _GEN_72 = nextBitValid ? outputMemBlock_14 : outputMemBlock_13;
  assign _GEN_73 = nextBitValid ? outputMemBlock_15 : outputMemBlock_14;
  assign _GEN_74 = nextBitValid ? _T_143 : outputPieceBits;
  assign _GEN_75 = nextBitValid ? _T_146 : outputBits;
  assign _T_148 = outputPieceBits == 5'h10;
  assign _T_151 = io_inputFinished & _T_79;
  assign _T_153 = outputPieceBits > 5'h0;
  assign _T_154 = _T_151 & _T_153;
  assign _T_155 = _T_148 | _T_154;
  assign _T_156 = {outputMemBlock_1,outputMemBlock_0};
  assign _T_157 = {outputMemBlock_3,outputMemBlock_2};
  assign _T_158 = {_T_157,_T_156};
  assign _T_159 = {outputMemBlock_5,outputMemBlock_4};
  assign _T_160 = {outputMemBlock_7,outputMemBlock_6};
  assign _T_161 = {_T_160,_T_159};
  assign _T_162 = {_T_161,_T_158};
  assign _T_163 = {outputMemBlock_9,outputMemBlock_8};
  assign _T_164 = {outputMemBlock_11,outputMemBlock_10};
  assign _T_165 = {_T_164,_T_163};
  assign _T_166 = {outputMemBlock_13,outputMemBlock_12};
  assign _T_167 = {outputMemBlock_15,outputMemBlock_14};
  assign _T_168 = {_T_167,_T_166};
  assign _T_169 = {_T_168,_T_165};
  assign _T_170 = {_T_169,_T_162};
  assign _T_175 = outputWriteAddr + 5'h1;
  assign _T_176 = _T_175[4:0];
  assign _GEN_76 = _T_148 ? 5'h0 : _GEN_74;
  assign _GEN_77 = _T_148 ? _T_176 : outputWriteAddr;
  assign _T_181 = outputReadingStarted == 1'h0;
  assign _T_188 = outputBits > 10'h0;
  assign _T_189 = _T_151 & _T_188;
  assign _T_190 = _T_122 | _T_189;
  assign _T_191 = _T_181 & _T_190;
  assign _GEN_78 = _T_191 ? 1'h1 : outputReadingStarted;
  assign _T_193 = io_outputMemBlockReady & outputReadingStarted;
  assign _T_195 = outputReadAddr != 5'h1f;
  assign _T_196 = _T_193 & _T_195;
  assign _T_198 = outputReadAddr + 5'h1;
  assign _T_199 = _T_198[4:0];
  assign _GEN_79 = _T_196 ? _T_199 : outputReadAddr;
  assign _T_203 = io_inputFinished == 1'h0;
  assign _T_204 = _T_79 & _T_203;
  assign _T_214 = outputReadingStarted & _T_190;
  assign _T_219 = outputBits == 10'h0;
  assign _T_220 = _T_151 & _T_219;
  assign _GEN_80 = io_outputMemFlushed ? 10'h0 : _GEN_75;
  assign _GEN_81 = io_outputMemFlushed ? 5'h0 : _GEN_76;
  assign _GEN_82 = io_outputMemFlushed ? 1'h0 : _GEN_78;
  assign _GEN_83 = io_outputMemFlushed ? 5'h0 : _GEN_77;
  assign _GEN_84 = io_outputMemFlushed ? 5'h0 : _GEN_79;
  assign io_inputMemConsumed = _T_204;
  assign io_outputMemBlock = outputBram_io_b_dout;
  assign io_outputMemBlockValid = _T_214;
  assign io_outputBits = outputBits;
  assign io_outputFinished = _T_220;
  assign inputBram_io_a_addr = io_inputMemIdx;
  assign inputBram_io_a_din = io_inputMemBlock;
  assign inputBram_io_a_wr = io_inputMemBlockValid;
  assign inputBram_io_b_addr = inputReadAddr;
  assign inputBram_clock = clock;
  assign outputBram_io_a_addr = outputWriteAddr;
  assign outputBram_io_a_din = _T_170;
  assign outputBram_io_a_wr = _T_155;
  assign outputBram_io_b_addr = outputReadAddr;
  assign outputBram_clock = clock;
  assign inputAdvance = _T_130;
  assign nextBitValid = inputAdvance;
  assign nextBit = inputMemBlock_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  inputMemBlock_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  inputMemBlock_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputMemBlock_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  inputMemBlock_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  inputMemBlock_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  inputMemBlock_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  inputMemBlock_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemBlock_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBlock_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  inputMemBlock_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputMemBlock_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  inputMemBlock_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  inputMemBlock_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  inputMemBlock_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  inputMemBlock_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  inputMemBlock_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  inputPieceBitsRemaining = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  inputBitsRemaining = _RAND_17[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  inputBlockLoaded = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  outputMemBlock_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  outputMemBlock_1 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  outputMemBlock_2 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  outputMemBlock_3 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  outputMemBlock_4 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  outputMemBlock_5 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  outputMemBlock_6 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  outputMemBlock_7 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  outputMemBlock_8 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  outputMemBlock_9 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  outputMemBlock_10 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  outputMemBlock_11 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  outputMemBlock_12 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  outputMemBlock_13 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  outputMemBlock_14 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  outputMemBlock_15 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  outputBits = _RAND_35[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  outputPieceBits = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  inputReadAddr = _RAND_37[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  inputPieceRead = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  outputWriteAddr = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  outputReadAddr = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  outputReadingStarted = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (inputAdvance) begin
      inputMemBlock_0 <= inputMemBlock_1;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_0 <= _T_102;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_1 <= inputMemBlock_2;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_1 <= _T_103;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_2 <= inputMemBlock_3;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_2 <= _T_104;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_3 <= inputMemBlock_4;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_3 <= _T_105;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_4 <= inputMemBlock_5;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_4 <= _T_106;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_5 <= inputMemBlock_6;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_5 <= _T_107;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_6 <= inputMemBlock_7;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_6 <= _T_108;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_7 <= inputMemBlock_8;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_7 <= _T_109;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_8 <= inputMemBlock_9;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_8 <= _T_110;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_9 <= inputMemBlock_10;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_9 <= _T_111;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_10 <= inputMemBlock_11;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_10 <= _T_112;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_11 <= inputMemBlock_12;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_11 <= _T_113;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_12 <= inputMemBlock_13;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_12 <= _T_114;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_13 <= inputMemBlock_14;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_13 <= _T_115;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_14 <= inputMemBlock_15;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_14 <= _T_116;
        end
      end
    end
    if (_T_90) begin
      if (!(_T_92)) begin
        inputMemBlock_15 <= _T_117;
      end
    end
    if (reset) begin
      inputPieceBitsRemaining <= 5'h0;
    end else begin
      inputPieceBitsRemaining <= _GEN_41[4:0];
    end
    if (reset) begin
      inputBitsRemaining <= 10'h0;
    end else begin
      if (inputAdvance) begin
        inputBitsRemaining <= _T_138;
      end else begin
        if (_T_76) begin
          inputBitsRemaining <= io_inputBits;
        end
      end
    end
    if (reset) begin
      inputBlockLoaded <= 1'h0;
    end else begin
      if (_T_80) begin
        inputBlockLoaded <= 1'h0;
      end else begin
        if (_T_76) begin
          inputBlockLoaded <= 1'h1;
        end
      end
    end
    if (nextBitValid) begin
      outputMemBlock_0 <= outputMemBlock_1;
    end
    if (nextBitValid) begin
      outputMemBlock_1 <= outputMemBlock_2;
    end
    if (nextBitValid) begin
      outputMemBlock_2 <= outputMemBlock_3;
    end
    if (nextBitValid) begin
      outputMemBlock_3 <= outputMemBlock_4;
    end
    if (nextBitValid) begin
      outputMemBlock_4 <= outputMemBlock_5;
    end
    if (nextBitValid) begin
      outputMemBlock_5 <= outputMemBlock_6;
    end
    if (nextBitValid) begin
      outputMemBlock_6 <= outputMemBlock_7;
    end
    if (nextBitValid) begin
      outputMemBlock_7 <= outputMemBlock_8;
    end
    if (nextBitValid) begin
      outputMemBlock_8 <= outputMemBlock_9;
    end
    if (nextBitValid) begin
      outputMemBlock_9 <= outputMemBlock_10;
    end
    if (nextBitValid) begin
      outputMemBlock_10 <= outputMemBlock_11;
    end
    if (nextBitValid) begin
      outputMemBlock_11 <= outputMemBlock_12;
    end
    if (nextBitValid) begin
      outputMemBlock_12 <= outputMemBlock_13;
    end
    if (nextBitValid) begin
      outputMemBlock_13 <= outputMemBlock_14;
    end
    if (nextBitValid) begin
      outputMemBlock_14 <= outputMemBlock_15;
    end
    if (nextBitValid) begin
      outputMemBlock_15 <= nextBit;
    end
    if (reset) begin
      outputBits <= 10'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputBits <= 10'h0;
      end else begin
        if (nextBitValid) begin
          outputBits <= _T_146;
        end
      end
    end
    if (reset) begin
      outputPieceBits <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputPieceBits <= 5'h0;
      end else begin
        if (_T_148) begin
          outputPieceBits <= 5'h0;
        end else begin
          if (nextBitValid) begin
            outputPieceBits <= _T_143;
          end
        end
      end
    end
    if (reset) begin
      inputReadAddr <= 5'h0;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputReadAddr <= _T_101;
        end
      end
    end
    if (reset) begin
      inputPieceRead <= 1'h0;
    end else begin
      if (_T_90) begin
        inputPieceRead <= _T_92;
      end
    end
    if (reset) begin
      outputWriteAddr <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputWriteAddr <= 5'h0;
      end else begin
        if (_T_148) begin
          outputWriteAddr <= _T_176;
        end
      end
    end
    if (reset) begin
      outputReadAddr <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputReadAddr <= 5'h0;
      end else begin
        if (_T_196) begin
          outputReadAddr <= _T_199;
        end
      end
    end
    if (reset) begin
      outputReadingStarted <= 1'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputReadingStarted <= 1'h0;
      end else begin
        if (_T_191) begin
          outputReadingStarted <= 1'h1;
        end
      end
    end
  end
endmodule
module StreamingCore(
  input         clock,
  input         reset,
  output [31:0] io_inputMemAddr,
  input         io_inputMemAddrConsumed,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output        io_inputMemBlockReady,
  output [31:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [15:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output        io_inputAddrsIgnore,
  output        io_inputBlocksFinished,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [15:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [15:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [31:0] inputBitsRemaining;
  reg [31:0] _RAND_2;
  reg  coreInputFinished;
  reg [31:0] _RAND_3;
  reg [31:0] outputBits;
  reg [31:0] _RAND_4;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_5;
  reg  outputLengthCommitted;
  reg [31:0] _RAND_6;
  reg [31:0] inputMemAddr;
  reg [31:0] _RAND_7;
  reg [31:0] inputMemBound;
  reg [31:0] _RAND_8;
  reg [31:0] outputMemAddr;
  reg [31:0] _RAND_9;
  reg [31:0] outputLenAddr;
  reg [31:0] _RAND_10;
  wire  _T_40;
  wire  _T_41;
  wire  _T_44;
  reg  initAddressAcked;
  reg [31:0] _RAND_11;
  wire  _GEN_0;
  wire  _T_48;
  wire [32:0] _T_50;
  wire [31:0] _T_51;
  wire [31:0] _GEN_1;
  wire  _T_52;
  wire  _T_53;
  wire  _T_54;
  wire  _T_55;
  wire  _T_57;
  wire  _T_59;
  wire  _T_60;
  wire  _T_61;
  wire  _T_62;
  wire  _T_64;
  wire [31:0] _T_66;
  wire  _T_68;
  wire [15:0] _T_69;
  wire [31:0] _T_70;
  wire [31:0] _GEN_2;
  wire  _T_72;
  wire [15:0] _T_73;
  wire [31:0] _T_74;
  wire [31:0] _GEN_3;
  wire  _T_76;
  wire [15:0] _T_77;
  wire [31:0] _T_78;
  wire [22:0] _T_79;
  wire [28:0] _T_81;
  wire [31:0] _GEN_44;
  wire [32:0] _T_82;
  wire [31:0] _T_83;
  wire [8:0] _T_84;
  wire  _T_86;
  wire [6:0] _T_89;
  wire [31:0] _GEN_45;
  wire [32:0] _T_90;
  wire [31:0] _T_91;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire  _T_93;
  wire [15:0] _T_94;
  wire [31:0] _T_95;
  wire [22:0] _T_96;
  wire [28:0] _T_98;
  wire [31:0] _GEN_46;
  wire [32:0] _T_99;
  wire [31:0] _T_100;
  wire [8:0] _T_101;
  wire  _T_103;
  wire [6:0] _T_106;
  wire [31:0] _GEN_47;
  wire [32:0] _T_107;
  wire [31:0] _T_108;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire  _T_110;
  wire [15:0] _T_111;
  wire [31:0] _T_112;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire  _T_114;
  wire [15:0] _T_115;
  wire [31:0] _T_116;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire  _T_118;
  wire [32:0] _T_122;
  wire [31:0] _T_123;
  wire  _GEN_12;
  wire  _GEN_13;
  wire [31:0] _GEN_14;
  wire [32:0] _T_129;
  wire [32:0] _T_130;
  wire [31:0] _T_131;
  wire [31:0] _T_133;
  wire [31:0] _GEN_15;
  wire [31:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [31:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [31:0] _GEN_23;
  wire [31:0] _GEN_24;
  wire [31:0] _GEN_25;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _T_138;
  wire  _GEN_30;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_12;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_13;
  wire  _GEN_31;
  wire [31:0] _T_145;
  wire  _T_147;
  wire  _T_149;
  wire  _T_150;
  wire  _T_151;
  wire  _T_152;
  wire  _T_153;
  wire  _GEN_32;
  wire  _T_159;
  wire [4:0] _GEN_33;
  wire [5:0] _T_162;
  wire [4:0] _T_163;
  wire [4:0] _GEN_34;
  wire [4:0] _GEN_35;
  wire [15:0] outputBitsBlock;
  wire  _T_166;
  wire [15:0] _T_167;
  wire  _T_169;
  wire [15:0] _T_170;
  wire [15:0] _T_172;
  wire [15:0] _T_173;
  wire [15:0] _T_174;
  wire  _T_175;
  wire  _T_179;
  wire [31:0] _GEN_48;
  wire [32:0] _T_183;
  wire [31:0] _T_184;
  wire  _GEN_36;
  wire [31:0] _GEN_37;
  wire [31:0] _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign _T_40 = io_inputAddrsIgnore == 1'h0;
  assign _T_41 = io_inputMemAddrConsumed & _T_40;
  assign _T_44 = reset == 1'h0;
  assign _GEN_0 = io_inputMemAddrConsumed ? 1'h1 : initAddressAcked;
  assign _T_48 = io_inputMemAddrConsumed & initDone;
  assign _T_50 = inputMemAddr + 32'h40;
  assign _T_51 = _T_50[31:0];
  assign _GEN_1 = _T_48 ? _T_51 : inputMemAddr;
  assign _T_52 = initAddressAcked & isInit;
  assign _T_53 = inputMemAddr == inputMemBound;
  assign _T_54 = _T_52 | _T_53;
  assign _T_55 = initDone & core_io_inputMemConsumed;
  assign _T_57 = inputBitsRemaining == 32'h0;
  assign _T_59 = _T_57 == 1'h0;
  assign _T_60 = _T_55 & _T_59;
  assign _T_61 = isInit | _T_60;
  assign _T_62 = io_inputMemBlockValid & initDone;
  assign _T_64 = inputBitsRemaining > 32'h200;
  assign _T_66 = _T_64 ? 32'h200 : inputBitsRemaining;
  assign _T_68 = io_inputMemIdx == 5'h0;
  assign _T_69 = inputMemAddr[31:16];
  assign _T_70 = {_T_69,io_inputMemBlock};
  assign _GEN_2 = _T_68 ? _T_70 : _GEN_1;
  assign _T_72 = io_inputMemIdx == 5'h1;
  assign _T_73 = inputMemAddr[15:0];
  assign _T_74 = {io_inputMemBlock,_T_73};
  assign _GEN_3 = _T_72 ? _T_74 : _GEN_2;
  assign _T_76 = io_inputMemIdx == 5'h4;
  assign _T_77 = inputBitsRemaining[31:16];
  assign _T_78 = {_T_77,io_inputMemBlock};
  assign _T_79 = _T_78[31:9];
  assign _T_81 = {_T_79,6'h0};
  assign _GEN_44 = {{3'd0}, _T_81};
  assign _T_82 = inputMemAddr + _GEN_44;
  assign _T_83 = _T_82[31:0];
  assign _T_84 = _T_78[8:0];
  assign _T_86 = _T_84 != 9'h0;
  assign _T_89 = _T_86 ? 7'h40 : 7'h0;
  assign _GEN_45 = {{25'd0}, _T_89};
  assign _T_90 = _T_83 + _GEN_45;
  assign _T_91 = _T_90[31:0];
  assign _GEN_4 = _T_76 ? _T_78 : inputBitsRemaining;
  assign _GEN_5 = _T_76 ? _T_91 : inputMemBound;
  assign _T_93 = io_inputMemIdx == 5'h5;
  assign _T_94 = inputBitsRemaining[15:0];
  assign _T_95 = {io_inputMemBlock,_T_94};
  assign _T_96 = _T_95[31:9];
  assign _T_98 = {_T_96,6'h0};
  assign _GEN_46 = {{3'd0}, _T_98};
  assign _T_99 = inputMemAddr + _GEN_46;
  assign _T_100 = _T_99[31:0];
  assign _T_101 = _T_95[8:0];
  assign _T_103 = _T_101 != 9'h0;
  assign _T_106 = _T_103 ? 7'h40 : 7'h0;
  assign _GEN_47 = {{25'd0}, _T_106};
  assign _T_107 = _T_100 + _GEN_47;
  assign _T_108 = _T_107[31:0];
  assign _GEN_6 = _T_93 ? _T_95 : _GEN_4;
  assign _GEN_7 = _T_93 ? _T_108 : _GEN_5;
  assign _T_110 = io_inputMemIdx == 5'h8;
  assign _T_111 = outputMemAddr[31:16];
  assign _T_112 = {_T_111,io_inputMemBlock};
  assign _GEN_8 = _T_110 ? _T_112 : outputMemAddr;
  assign _GEN_9 = _T_110 ? _T_112 : outputLenAddr;
  assign _T_114 = io_inputMemIdx == 5'h9;
  assign _T_115 = outputMemAddr[15:0];
  assign _T_116 = {io_inputMemBlock,_T_115};
  assign _GEN_10 = _T_114 ? _T_116 : _GEN_8;
  assign _GEN_11 = _T_114 ? _T_116 : _GEN_9;
  assign _T_118 = io_inputMemIdx == 5'h1f;
  assign _T_122 = outputMemAddr + 32'h40;
  assign _T_123 = _T_122[31:0];
  assign _GEN_12 = _T_118 ? 1'h0 : isInit;
  assign _GEN_13 = _T_118 ? 1'h1 : initDone;
  assign _GEN_14 = _T_118 ? _T_123 : _GEN_10;
  assign _T_129 = inputBitsRemaining - 32'h200;
  assign _T_130 = $unsigned(_T_129);
  assign _T_131 = _T_130[31:0];
  assign _T_133 = _T_64 ? _T_131 : 32'h0;
  assign _GEN_15 = _T_118 ? _T_133 : inputBitsRemaining;
  assign _GEN_16 = isInit ? _GEN_3 : _GEN_1;
  assign _GEN_17 = isInit ? _GEN_6 : _GEN_15;
  assign _GEN_18 = isInit ? _GEN_7 : inputMemBound;
  assign _GEN_19 = isInit ? _GEN_14 : outputMemAddr;
  assign _GEN_20 = isInit ? _GEN_11 : outputLenAddr;
  assign _GEN_21 = isInit ? _GEN_12 : isInit;
  assign _GEN_22 = isInit ? _GEN_13 : initDone;
  assign _GEN_23 = io_inputMemBlockValid ? _GEN_16 : _GEN_1;
  assign _GEN_24 = io_inputMemBlockValid ? _GEN_17 : inputBitsRemaining;
  assign _GEN_25 = io_inputMemBlockValid ? _GEN_18 : inputMemBound;
  assign _GEN_26 = io_inputMemBlockValid ? _GEN_19 : outputMemAddr;
  assign _GEN_27 = io_inputMemBlockValid ? _GEN_20 : outputLenAddr;
  assign _GEN_28 = io_inputMemBlockValid ? _GEN_21 : isInit;
  assign _GEN_29 = io_inputMemBlockValid ? _GEN_22 : initDone;
  assign _T_138 = core_io_inputMemConsumed & _T_57;
  assign _GEN_30 = _T_138 ? 1'h1 : coreInputFinished;
  assign _GEN_31 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_145 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_147 = outputAddressAccepted == 1'h0;
  assign _T_149 = outputLengthCommitted == 1'h0;
  assign _T_150 = core_io_outputFinished & _T_149;
  assign _T_151 = core_io_outputMemBlockValid | _T_150;
  assign _T_152 = _T_147 & _T_151;
  assign _T_153 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_32 = _T_153 ? 1'h1 : outputAddressAccepted;
  assign _T_159 = outputBlockCounter == 5'h1f;
  assign _GEN_33 = io_outputMemBlockReady ? 5'h0 : outputBlockCounter;
  assign _T_162 = outputBlockCounter + 5'h1;
  assign _T_163 = _T_162[4:0];
  assign _GEN_34 = _T_159 ? _GEN_33 : _T_163;
  assign _GEN_35 = outputAddressAcceptedNext ? _GEN_34 : outputBlockCounter;
  assign _T_166 = outputBlockCounter == 5'h0;
  assign _T_167 = outputBits[15:0];
  assign _T_169 = outputBlockCounter == 5'h1;
  assign _T_170 = outputBits[31:16];
  assign _T_172 = _T_169 ? _T_170 : 16'h0;
  assign _T_173 = _T_166 ? _T_167 : _T_172;
  assign _T_174 = core_io_outputFinished ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_175 = outputAddressAcceptedNext & io_outputMemBlockReady;
  assign _T_179 = _T_175 & _T_159;
  assign _GEN_48 = {{22'd0}, core_io_outputBits};
  assign _T_183 = outputBits + _GEN_48;
  assign _T_184 = _T_183[31:0];
  assign _GEN_36 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _GEN_37 = core_io_outputFinished ? outputBits : _T_184;
  assign _GEN_38 = core_io_outputFinished ? _GEN_26 : _T_123;
  assign _GEN_39 = _T_179 ? 1'h0 : _GEN_32;
  assign _GEN_40 = _T_179 ? 1'h0 : _GEN_31;
  assign _GEN_41 = _T_179 ? _GEN_36 : outputLengthCommitted;
  assign _GEN_42 = _T_179 ? _GEN_37 : outputBits;
  assign _GEN_43 = _T_179 ? _GEN_38 : _GEN_26;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemBlockReady = _T_61;
  assign io_outputMemAddr = _T_145;
  assign io_outputMemAddrValid = _T_152;
  assign io_outputMemBlock = _T_174;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_inputAddrsIgnore = _T_54;
  assign io_inputBlocksFinished = _T_57;
  assign io_outputFinished = outputLengthCommitted;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_62;
  assign core_io_inputBits = _T_66[9:0];
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_io_outputMemFlushed = _T_175;
  assign core_clock = clock;
  assign core_reset = reset;
  assign outputBitsBlock = _T_173;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputBitsRemaining = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  coreInputFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  outputBits = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputBlockCounter = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputLengthCommitted = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemAddr = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBound = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  outputMemAddr = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  outputLenAddr = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  initAddressAcked = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  outputAddressAccepted = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  outputAddressAcceptedNext = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_118) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_118) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 32'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_93) begin
            inputBitsRemaining <= _T_95;
          end else begin
            if (_T_76) begin
              inputBitsRemaining <= _T_78;
            end
          end
        end else begin
          if (_T_118) begin
            if (_T_64) begin
              inputBitsRemaining <= _T_131;
            end else begin
              inputBitsRemaining <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_138) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 32'h0;
    end else begin
      if (_T_179) begin
        if (!(core_io_outputFinished)) begin
          outputBits <= _T_184;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_159) begin
          if (io_outputMemBlockReady) begin
            outputBlockCounter <= 5'h0;
          end
        end else begin
          outputBlockCounter <= _T_163;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_179) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 32'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_72) begin
            inputMemAddr <= _T_74;
          end else begin
            if (_T_68) begin
              inputMemAddr <= _T_70;
            end else begin
              if (_T_48) begin
                inputMemAddr <= _T_51;
              end
            end
          end
        end else begin
          if (_T_48) begin
            inputMemAddr <= _T_51;
          end
        end
      end else begin
        if (_T_48) begin
          inputMemAddr <= _T_51;
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_93) begin
          inputMemBound <= _T_108;
        end else begin
          if (_T_76) begin
            inputMemBound <= _T_91;
          end
        end
      end
    end
    if (_T_179) begin
      if (core_io_outputFinished) begin
        if (io_inputMemBlockValid) begin
          if (isInit) begin
            if (_T_118) begin
              outputMemAddr <= _T_123;
            end else begin
              if (_T_114) begin
                outputMemAddr <= _T_116;
              end else begin
                if (_T_110) begin
                  outputMemAddr <= _T_112;
                end
              end
            end
          end
        end
      end else begin
        outputMemAddr <= _T_123;
      end
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_118) begin
            outputMemAddr <= _T_123;
          end else begin
            if (_T_114) begin
              outputMemAddr <= _T_116;
            end else begin
              if (_T_110) begin
                outputMemAddr <= _T_112;
              end
            end
          end
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_114) begin
          outputLenAddr <= _T_116;
        end else begin
          if (_T_110) begin
            outputLenAddr <= _T_112;
          end
        end
      end
    end
    if (reset) begin
      initAddressAcked <= 1'h0;
    end else begin
      if (io_inputMemAddrConsumed) begin
        initAddressAcked <= 1'h1;
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_179) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_153) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_179) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41 & _T_44) begin
          $fwrite(32'h80000002,"input address 0x%h accepted for core 0\n",io_inputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_153 & _T_44) begin
          $fwrite(32'h80000002,"output address 0x%h accepted for core 0\n",io_outputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module StreamingCore_1(
  input         clock,
  input         reset,
  output [31:0] io_inputMemAddr,
  input         io_inputMemAddrConsumed,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output        io_inputMemBlockReady,
  output [31:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [15:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output        io_inputAddrsIgnore,
  output        io_inputBlocksFinished,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [15:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [15:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [31:0] inputBitsRemaining;
  reg [31:0] _RAND_2;
  reg  coreInputFinished;
  reg [31:0] _RAND_3;
  reg [31:0] outputBits;
  reg [31:0] _RAND_4;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_5;
  reg  outputLengthCommitted;
  reg [31:0] _RAND_6;
  reg [31:0] inputMemAddr;
  reg [31:0] _RAND_7;
  reg [31:0] inputMemBound;
  reg [31:0] _RAND_8;
  reg [31:0] outputMemAddr;
  reg [31:0] _RAND_9;
  reg [31:0] outputLenAddr;
  reg [31:0] _RAND_10;
  wire  _T_40;
  wire  _T_41;
  wire  _T_44;
  reg  initAddressAcked;
  reg [31:0] _RAND_11;
  wire  _GEN_0;
  wire  _T_48;
  wire [32:0] _T_50;
  wire [31:0] _T_51;
  wire [31:0] _GEN_1;
  wire  _T_52;
  wire  _T_53;
  wire  _T_54;
  wire  _T_55;
  wire  _T_57;
  wire  _T_59;
  wire  _T_60;
  wire  _T_61;
  wire  _T_62;
  wire  _T_64;
  wire [31:0] _T_66;
  wire  _T_68;
  wire [15:0] _T_69;
  wire [31:0] _T_70;
  wire [31:0] _GEN_2;
  wire  _T_72;
  wire [15:0] _T_73;
  wire [31:0] _T_74;
  wire [31:0] _GEN_3;
  wire  _T_76;
  wire [15:0] _T_77;
  wire [31:0] _T_78;
  wire [22:0] _T_79;
  wire [28:0] _T_81;
  wire [31:0] _GEN_44;
  wire [32:0] _T_82;
  wire [31:0] _T_83;
  wire [8:0] _T_84;
  wire  _T_86;
  wire [6:0] _T_89;
  wire [31:0] _GEN_45;
  wire [32:0] _T_90;
  wire [31:0] _T_91;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire  _T_93;
  wire [15:0] _T_94;
  wire [31:0] _T_95;
  wire [22:0] _T_96;
  wire [28:0] _T_98;
  wire [31:0] _GEN_46;
  wire [32:0] _T_99;
  wire [31:0] _T_100;
  wire [8:0] _T_101;
  wire  _T_103;
  wire [6:0] _T_106;
  wire [31:0] _GEN_47;
  wire [32:0] _T_107;
  wire [31:0] _T_108;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire  _T_110;
  wire [15:0] _T_111;
  wire [31:0] _T_112;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire  _T_114;
  wire [15:0] _T_115;
  wire [31:0] _T_116;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire  _T_118;
  wire [32:0] _T_122;
  wire [31:0] _T_123;
  wire  _GEN_12;
  wire  _GEN_13;
  wire [31:0] _GEN_14;
  wire [32:0] _T_129;
  wire [32:0] _T_130;
  wire [31:0] _T_131;
  wire [31:0] _T_133;
  wire [31:0] _GEN_15;
  wire [31:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [31:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [31:0] _GEN_23;
  wire [31:0] _GEN_24;
  wire [31:0] _GEN_25;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _T_138;
  wire  _GEN_30;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_12;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_13;
  wire  _GEN_31;
  wire [31:0] _T_145;
  wire  _T_147;
  wire  _T_149;
  wire  _T_150;
  wire  _T_151;
  wire  _T_152;
  wire  _T_153;
  wire  _GEN_32;
  wire  _T_159;
  wire [4:0] _GEN_33;
  wire [5:0] _T_162;
  wire [4:0] _T_163;
  wire [4:0] _GEN_34;
  wire [4:0] _GEN_35;
  wire [15:0] outputBitsBlock;
  wire  _T_166;
  wire [15:0] _T_167;
  wire  _T_169;
  wire [15:0] _T_170;
  wire [15:0] _T_172;
  wire [15:0] _T_173;
  wire [15:0] _T_174;
  wire  _T_175;
  wire  _T_179;
  wire [31:0] _GEN_48;
  wire [32:0] _T_183;
  wire [31:0] _T_184;
  wire  _GEN_36;
  wire [31:0] _GEN_37;
  wire [31:0] _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign _T_40 = io_inputAddrsIgnore == 1'h0;
  assign _T_41 = io_inputMemAddrConsumed & _T_40;
  assign _T_44 = reset == 1'h0;
  assign _GEN_0 = io_inputMemAddrConsumed ? 1'h1 : initAddressAcked;
  assign _T_48 = io_inputMemAddrConsumed & initDone;
  assign _T_50 = inputMemAddr + 32'h40;
  assign _T_51 = _T_50[31:0];
  assign _GEN_1 = _T_48 ? _T_51 : inputMemAddr;
  assign _T_52 = initAddressAcked & isInit;
  assign _T_53 = inputMemAddr == inputMemBound;
  assign _T_54 = _T_52 | _T_53;
  assign _T_55 = initDone & core_io_inputMemConsumed;
  assign _T_57 = inputBitsRemaining == 32'h0;
  assign _T_59 = _T_57 == 1'h0;
  assign _T_60 = _T_55 & _T_59;
  assign _T_61 = isInit | _T_60;
  assign _T_62 = io_inputMemBlockValid & initDone;
  assign _T_64 = inputBitsRemaining > 32'h200;
  assign _T_66 = _T_64 ? 32'h200 : inputBitsRemaining;
  assign _T_68 = io_inputMemIdx == 5'h0;
  assign _T_69 = inputMemAddr[31:16];
  assign _T_70 = {_T_69,io_inputMemBlock};
  assign _GEN_2 = _T_68 ? _T_70 : _GEN_1;
  assign _T_72 = io_inputMemIdx == 5'h1;
  assign _T_73 = inputMemAddr[15:0];
  assign _T_74 = {io_inputMemBlock,_T_73};
  assign _GEN_3 = _T_72 ? _T_74 : _GEN_2;
  assign _T_76 = io_inputMemIdx == 5'h4;
  assign _T_77 = inputBitsRemaining[31:16];
  assign _T_78 = {_T_77,io_inputMemBlock};
  assign _T_79 = _T_78[31:9];
  assign _T_81 = {_T_79,6'h0};
  assign _GEN_44 = {{3'd0}, _T_81};
  assign _T_82 = inputMemAddr + _GEN_44;
  assign _T_83 = _T_82[31:0];
  assign _T_84 = _T_78[8:0];
  assign _T_86 = _T_84 != 9'h0;
  assign _T_89 = _T_86 ? 7'h40 : 7'h0;
  assign _GEN_45 = {{25'd0}, _T_89};
  assign _T_90 = _T_83 + _GEN_45;
  assign _T_91 = _T_90[31:0];
  assign _GEN_4 = _T_76 ? _T_78 : inputBitsRemaining;
  assign _GEN_5 = _T_76 ? _T_91 : inputMemBound;
  assign _T_93 = io_inputMemIdx == 5'h5;
  assign _T_94 = inputBitsRemaining[15:0];
  assign _T_95 = {io_inputMemBlock,_T_94};
  assign _T_96 = _T_95[31:9];
  assign _T_98 = {_T_96,6'h0};
  assign _GEN_46 = {{3'd0}, _T_98};
  assign _T_99 = inputMemAddr + _GEN_46;
  assign _T_100 = _T_99[31:0];
  assign _T_101 = _T_95[8:0];
  assign _T_103 = _T_101 != 9'h0;
  assign _T_106 = _T_103 ? 7'h40 : 7'h0;
  assign _GEN_47 = {{25'd0}, _T_106};
  assign _T_107 = _T_100 + _GEN_47;
  assign _T_108 = _T_107[31:0];
  assign _GEN_6 = _T_93 ? _T_95 : _GEN_4;
  assign _GEN_7 = _T_93 ? _T_108 : _GEN_5;
  assign _T_110 = io_inputMemIdx == 5'h8;
  assign _T_111 = outputMemAddr[31:16];
  assign _T_112 = {_T_111,io_inputMemBlock};
  assign _GEN_8 = _T_110 ? _T_112 : outputMemAddr;
  assign _GEN_9 = _T_110 ? _T_112 : outputLenAddr;
  assign _T_114 = io_inputMemIdx == 5'h9;
  assign _T_115 = outputMemAddr[15:0];
  assign _T_116 = {io_inputMemBlock,_T_115};
  assign _GEN_10 = _T_114 ? _T_116 : _GEN_8;
  assign _GEN_11 = _T_114 ? _T_116 : _GEN_9;
  assign _T_118 = io_inputMemIdx == 5'h1f;
  assign _T_122 = outputMemAddr + 32'h40;
  assign _T_123 = _T_122[31:0];
  assign _GEN_12 = _T_118 ? 1'h0 : isInit;
  assign _GEN_13 = _T_118 ? 1'h1 : initDone;
  assign _GEN_14 = _T_118 ? _T_123 : _GEN_10;
  assign _T_129 = inputBitsRemaining - 32'h200;
  assign _T_130 = $unsigned(_T_129);
  assign _T_131 = _T_130[31:0];
  assign _T_133 = _T_64 ? _T_131 : 32'h0;
  assign _GEN_15 = _T_118 ? _T_133 : inputBitsRemaining;
  assign _GEN_16 = isInit ? _GEN_3 : _GEN_1;
  assign _GEN_17 = isInit ? _GEN_6 : _GEN_15;
  assign _GEN_18 = isInit ? _GEN_7 : inputMemBound;
  assign _GEN_19 = isInit ? _GEN_14 : outputMemAddr;
  assign _GEN_20 = isInit ? _GEN_11 : outputLenAddr;
  assign _GEN_21 = isInit ? _GEN_12 : isInit;
  assign _GEN_22 = isInit ? _GEN_13 : initDone;
  assign _GEN_23 = io_inputMemBlockValid ? _GEN_16 : _GEN_1;
  assign _GEN_24 = io_inputMemBlockValid ? _GEN_17 : inputBitsRemaining;
  assign _GEN_25 = io_inputMemBlockValid ? _GEN_18 : inputMemBound;
  assign _GEN_26 = io_inputMemBlockValid ? _GEN_19 : outputMemAddr;
  assign _GEN_27 = io_inputMemBlockValid ? _GEN_20 : outputLenAddr;
  assign _GEN_28 = io_inputMemBlockValid ? _GEN_21 : isInit;
  assign _GEN_29 = io_inputMemBlockValid ? _GEN_22 : initDone;
  assign _T_138 = core_io_inputMemConsumed & _T_57;
  assign _GEN_30 = _T_138 ? 1'h1 : coreInputFinished;
  assign _GEN_31 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_145 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_147 = outputAddressAccepted == 1'h0;
  assign _T_149 = outputLengthCommitted == 1'h0;
  assign _T_150 = core_io_outputFinished & _T_149;
  assign _T_151 = core_io_outputMemBlockValid | _T_150;
  assign _T_152 = _T_147 & _T_151;
  assign _T_153 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_32 = _T_153 ? 1'h1 : outputAddressAccepted;
  assign _T_159 = outputBlockCounter == 5'h1f;
  assign _GEN_33 = io_outputMemBlockReady ? 5'h0 : outputBlockCounter;
  assign _T_162 = outputBlockCounter + 5'h1;
  assign _T_163 = _T_162[4:0];
  assign _GEN_34 = _T_159 ? _GEN_33 : _T_163;
  assign _GEN_35 = outputAddressAcceptedNext ? _GEN_34 : outputBlockCounter;
  assign _T_166 = outputBlockCounter == 5'h0;
  assign _T_167 = outputBits[15:0];
  assign _T_169 = outputBlockCounter == 5'h1;
  assign _T_170 = outputBits[31:16];
  assign _T_172 = _T_169 ? _T_170 : 16'h0;
  assign _T_173 = _T_166 ? _T_167 : _T_172;
  assign _T_174 = core_io_outputFinished ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_175 = outputAddressAcceptedNext & io_outputMemBlockReady;
  assign _T_179 = _T_175 & _T_159;
  assign _GEN_48 = {{22'd0}, core_io_outputBits};
  assign _T_183 = outputBits + _GEN_48;
  assign _T_184 = _T_183[31:0];
  assign _GEN_36 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _GEN_37 = core_io_outputFinished ? outputBits : _T_184;
  assign _GEN_38 = core_io_outputFinished ? _GEN_26 : _T_123;
  assign _GEN_39 = _T_179 ? 1'h0 : _GEN_32;
  assign _GEN_40 = _T_179 ? 1'h0 : _GEN_31;
  assign _GEN_41 = _T_179 ? _GEN_36 : outputLengthCommitted;
  assign _GEN_42 = _T_179 ? _GEN_37 : outputBits;
  assign _GEN_43 = _T_179 ? _GEN_38 : _GEN_26;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemBlockReady = _T_61;
  assign io_outputMemAddr = _T_145;
  assign io_outputMemAddrValid = _T_152;
  assign io_outputMemBlock = _T_174;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_inputAddrsIgnore = _T_54;
  assign io_inputBlocksFinished = _T_57;
  assign io_outputFinished = outputLengthCommitted;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_62;
  assign core_io_inputBits = _T_66[9:0];
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_io_outputMemFlushed = _T_175;
  assign core_clock = clock;
  assign core_reset = reset;
  assign outputBitsBlock = _T_173;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputBitsRemaining = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  coreInputFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  outputBits = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputBlockCounter = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputLengthCommitted = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemAddr = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBound = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  outputMemAddr = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  outputLenAddr = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  initAddressAcked = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  outputAddressAccepted = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  outputAddressAcceptedNext = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_118) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_118) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 32'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_93) begin
            inputBitsRemaining <= _T_95;
          end else begin
            if (_T_76) begin
              inputBitsRemaining <= _T_78;
            end
          end
        end else begin
          if (_T_118) begin
            if (_T_64) begin
              inputBitsRemaining <= _T_131;
            end else begin
              inputBitsRemaining <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_138) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 32'h0;
    end else begin
      if (_T_179) begin
        if (!(core_io_outputFinished)) begin
          outputBits <= _T_184;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_159) begin
          if (io_outputMemBlockReady) begin
            outputBlockCounter <= 5'h0;
          end
        end else begin
          outputBlockCounter <= _T_163;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_179) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 32'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_72) begin
            inputMemAddr <= _T_74;
          end else begin
            if (_T_68) begin
              inputMemAddr <= _T_70;
            end else begin
              if (_T_48) begin
                inputMemAddr <= _T_51;
              end
            end
          end
        end else begin
          if (_T_48) begin
            inputMemAddr <= _T_51;
          end
        end
      end else begin
        if (_T_48) begin
          inputMemAddr <= _T_51;
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_93) begin
          inputMemBound <= _T_108;
        end else begin
          if (_T_76) begin
            inputMemBound <= _T_91;
          end
        end
      end
    end
    if (_T_179) begin
      if (core_io_outputFinished) begin
        if (io_inputMemBlockValid) begin
          if (isInit) begin
            if (_T_118) begin
              outputMemAddr <= _T_123;
            end else begin
              if (_T_114) begin
                outputMemAddr <= _T_116;
              end else begin
                if (_T_110) begin
                  outputMemAddr <= _T_112;
                end
              end
            end
          end
        end
      end else begin
        outputMemAddr <= _T_123;
      end
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_118) begin
            outputMemAddr <= _T_123;
          end else begin
            if (_T_114) begin
              outputMemAddr <= _T_116;
            end else begin
              if (_T_110) begin
                outputMemAddr <= _T_112;
              end
            end
          end
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_114) begin
          outputLenAddr <= _T_116;
        end else begin
          if (_T_110) begin
            outputLenAddr <= _T_112;
          end
        end
      end
    end
    if (reset) begin
      initAddressAcked <= 1'h0;
    end else begin
      if (io_inputMemAddrConsumed) begin
        initAddressAcked <= 1'h1;
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_179) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_153) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_179) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41 & _T_44) begin
          $fwrite(32'h80000002,"input address 0x%h accepted for core 1\n",io_inputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_153 & _T_44) begin
          $fwrite(32'h80000002,"output address 0x%h accepted for core 1\n",io_outputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module StreamingWrapper(
  input          clock,
  input          reset,
  output [63:0]  io_inputMemAddrs_0,
  output [63:0]  io_inputMemAddrs_1,
  output         io_inputMemAddrValids_0,
  output         io_inputMemAddrValids_1,
  input          io_inputMemAddrReadys_0,
  input          io_inputMemAddrReadys_1,
  input  [511:0] io_inputMemBlocks_0,
  input  [511:0] io_inputMemBlocks_1,
  input          io_inputMemBlockValids_0,
  input          io_inputMemBlockValids_1,
  output         io_inputMemBlockReadys_0,
  output         io_inputMemBlockReadys_1,
  output [63:0]  io_outputMemAddrs_0,
  output [63:0]  io_outputMemAddrs_1,
  output         io_outputMemAddrValids_0,
  output         io_outputMemAddrValids_1,
  input          io_outputMemAddrReadys_0,
  input          io_outputMemAddrReadys_1,
  output [511:0] io_outputMemBlocks_0,
  output [511:0] io_outputMemBlocks_1,
  output         io_outputMemBlockValids_0,
  output         io_outputMemBlockValids_1,
  input          io_outputMemBlockReadys_0,
  input          io_outputMemBlockReadys_1,
  output         io_finished
);
  wire  StreamingCore_clock;
  wire  StreamingCore_reset;
  wire [31:0] StreamingCore_io_inputMemAddr;
  wire  StreamingCore_io_inputMemAddrConsumed;
  wire [15:0] StreamingCore_io_inputMemBlock;
  wire [4:0] StreamingCore_io_inputMemIdx;
  wire  StreamingCore_io_inputMemBlockValid;
  wire  StreamingCore_io_inputMemBlockReady;
  wire [31:0] StreamingCore_io_outputMemAddr;
  wire  StreamingCore_io_outputMemAddrValid;
  wire  StreamingCore_io_outputMemAddrReady;
  wire [15:0] StreamingCore_io_outputMemBlock;
  wire [4:0] StreamingCore_io_outputMemIdx;
  wire  StreamingCore_io_outputMemBlockValid;
  wire  StreamingCore_io_outputMemBlockReady;
  wire  StreamingCore_io_inputAddrsIgnore;
  wire  StreamingCore_io_inputBlocksFinished;
  wire  StreamingCore_io_outputFinished;
  wire  StreamingCore_1_clock;
  wire  StreamingCore_1_reset;
  wire [31:0] StreamingCore_1_io_inputMemAddr;
  wire  StreamingCore_1_io_inputMemAddrConsumed;
  wire [15:0] StreamingCore_1_io_inputMemBlock;
  wire [4:0] StreamingCore_1_io_inputMemIdx;
  wire  StreamingCore_1_io_inputMemBlockValid;
  wire  StreamingCore_1_io_inputMemBlockReady;
  wire [31:0] StreamingCore_1_io_outputMemAddr;
  wire  StreamingCore_1_io_outputMemAddrValid;
  wire  StreamingCore_1_io_outputMemAddrReady;
  wire [15:0] StreamingCore_1_io_outputMemBlock;
  wire [4:0] StreamingCore_1_io_outputMemIdx;
  wire  StreamingCore_1_io_outputMemBlockValid;
  wire  StreamingCore_1_io_outputMemBlockReady;
  wire  StreamingCore_1_io_inputAddrsIgnore;
  wire  StreamingCore_1_io_inputBlocksFinished;
  wire  StreamingCore_1_io_outputFinished;
  wire [31:0] cores_0_inputMemAddr;
  wire  cores_0_inputMemAddrConsumed;
  wire [15:0] cores_0_inputMemBlock;
  wire [4:0] cores_0_inputMemIdx;
  wire  cores_0_inputMemBlockValid;
  wire  cores_0_inputMemBlockReady;
  wire [31:0] cores_0_outputMemAddr;
  wire  cores_0_outputMemAddrValid;
  wire  cores_0_outputMemAddrReady;
  wire [15:0] cores_0_outputMemBlock;
  wire [4:0] cores_0_outputMemIdx;
  wire  cores_0_outputMemBlockValid;
  wire  cores_0_outputMemBlockReady;
  wire  cores_0_inputAddrsIgnore;
  wire  cores_0_inputBlocksFinished;
  wire  cores_0_outputFinished;
  wire [31:0] cores_1_inputMemAddr;
  wire  cores_1_inputMemAddrConsumed;
  wire [15:0] cores_1_inputMemBlock;
  wire [4:0] cores_1_inputMemIdx;
  wire  cores_1_inputMemBlockValid;
  wire  cores_1_inputMemBlockReady;
  wire [31:0] cores_1_outputMemAddr;
  wire  cores_1_outputMemAddrValid;
  wire  cores_1_outputMemAddrReady;
  wire [15:0] cores_1_outputMemBlock;
  wire [4:0] cores_1_outputMemIdx;
  wire  cores_1_outputMemBlockValid;
  wire  cores_1_outputMemBlockReady;
  wire  cores_1_inputAddrsIgnore;
  wire  cores_1_inputBlocksFinished;
  wire  cores_1_outputFinished;
  reg  _T_239;
  reg [31:0] _RAND_0;
  reg  _T_242;
  reg [31:0] _RAND_1;
  reg  _T_245;
  reg [31:0] _RAND_2;
  reg  _T_248;
  reg [31:0] _RAND_3;
  reg  _T_251;
  reg [31:0] _RAND_4;
  reg  _T_254;
  reg [31:0] _RAND_5;
  reg [63:0] _T_256;
  reg [63:0] _RAND_6;
  reg  _T_258;
  reg [31:0] _RAND_7;
  reg  _T_260;
  reg [31:0] _RAND_8;
  reg  _T_262;
  reg [31:0] _RAND_9;
  wire [63:0] _T_265_0;
  wire  _T_271_0;
  wire  _T_277_0;
  wire  _T_283_0;
  reg [63:0] _T_288;
  reg [63:0] _RAND_10;
  reg  _T_290;
  reg [31:0] _RAND_11;
  reg  _T_292;
  reg [31:0] _RAND_12;
  reg  _T_294;
  reg [31:0] _RAND_13;
  wire [63:0] _T_297_0;
  wire  _T_303_0;
  wire  _T_309_0;
  wire  _T_315_0;
  reg [63:0] _T_320;
  reg [63:0] _RAND_14;
  reg  _T_322;
  reg [31:0] _RAND_15;
  reg  _T_324;
  reg [31:0] _RAND_16;
  reg [15:0] _T_326;
  reg [31:0] _RAND_17;
  reg [4:0] _T_328;
  reg [31:0] _RAND_18;
  reg  _T_330;
  reg [31:0] _RAND_19;
  reg [63:0] _T_332;
  reg [63:0] _RAND_20;
  reg  _T_334;
  reg [31:0] _RAND_21;
  reg  _T_336;
  reg [31:0] _RAND_22;
  reg [15:0] _T_338;
  reg [31:0] _RAND_23;
  reg [4:0] _T_340;
  reg [31:0] _RAND_24;
  reg  _T_342;
  reg [31:0] _RAND_25;
  reg  _T_345;
  reg [31:0] _RAND_26;
  wire  _T_347;
  wire [1:0] _T_349;
  wire  _T_350;
  wire  _GEN_4;
  reg  _T_353;
  reg [31:0] _RAND_27;
  wire  _T_358;
  wire  _T_359;
  wire  _T_361;
  wire  _T_363;
  wire [1:0] _T_366;
  wire  _T_367;
  wire  _T_368;
  wire [1:0] _T_372;
  wire  _T_373;
  wire  _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _T_381;
  wire  _T_382;
  reg  _T_385;
  reg [31:0] _RAND_28;
  wire  _T_387;
  wire [1:0] _T_389;
  wire  _T_390;
  wire  _GEN_11;
  reg [15:0] _T_464_0_0;
  reg [31:0] _RAND_29;
  reg [15:0] _T_464_0_1;
  reg [31:0] _RAND_30;
  reg [15:0] _T_464_0_2;
  reg [31:0] _RAND_31;
  reg [15:0] _T_464_0_3;
  reg [31:0] _RAND_32;
  reg [15:0] _T_464_0_4;
  reg [31:0] _RAND_33;
  reg [15:0] _T_464_0_5;
  reg [31:0] _RAND_34;
  reg [15:0] _T_464_0_6;
  reg [31:0] _RAND_35;
  reg [15:0] _T_464_0_7;
  reg [31:0] _RAND_36;
  reg [15:0] _T_464_0_8;
  reg [31:0] _RAND_37;
  reg [15:0] _T_464_0_9;
  reg [31:0] _RAND_38;
  reg [15:0] _T_464_0_10;
  reg [31:0] _RAND_39;
  reg [15:0] _T_464_0_11;
  reg [31:0] _RAND_40;
  reg [15:0] _T_464_0_12;
  reg [31:0] _RAND_41;
  reg [15:0] _T_464_0_13;
  reg [31:0] _RAND_42;
  reg [15:0] _T_464_0_14;
  reg [31:0] _RAND_43;
  reg [15:0] _T_464_0_15;
  reg [31:0] _RAND_44;
  reg [15:0] _T_464_0_16;
  reg [31:0] _RAND_45;
  reg [15:0] _T_464_0_17;
  reg [31:0] _RAND_46;
  reg [15:0] _T_464_0_18;
  reg [31:0] _RAND_47;
  reg [15:0] _T_464_0_19;
  reg [31:0] _RAND_48;
  reg [15:0] _T_464_0_20;
  reg [31:0] _RAND_49;
  reg [15:0] _T_464_0_21;
  reg [31:0] _RAND_50;
  reg [15:0] _T_464_0_22;
  reg [31:0] _RAND_51;
  reg [15:0] _T_464_0_23;
  reg [31:0] _RAND_52;
  reg [15:0] _T_464_0_24;
  reg [31:0] _RAND_53;
  reg [15:0] _T_464_0_25;
  reg [31:0] _RAND_54;
  reg [15:0] _T_464_0_26;
  reg [31:0] _RAND_55;
  reg [15:0] _T_464_0_27;
  reg [31:0] _RAND_56;
  reg [15:0] _T_464_0_28;
  reg [31:0] _RAND_57;
  reg [15:0] _T_464_0_29;
  reg [31:0] _RAND_58;
  reg [15:0] _T_464_0_30;
  reg [31:0] _RAND_59;
  reg [15:0] _T_464_0_31;
  reg [31:0] _RAND_60;
  reg [4:0] _T_683_0;
  reg [31:0] _RAND_61;
  reg  _T_704_0;
  reg [31:0] _RAND_62;
  reg  _T_714;
  reg [31:0] _RAND_63;
  wire  _T_720;
  wire  _T_721;
  wire  _T_722;
  wire  _T_725;
  wire  _T_726;
  wire [15:0] _T_830;
  wire [15:0] _T_934;
  wire [15:0] _T_1038;
  wire [15:0] _T_1142;
  wire [15:0] _T_1246;
  wire [15:0] _T_1350;
  wire [15:0] _T_1454;
  wire [15:0] _T_1558;
  wire [15:0] _T_1662;
  wire [15:0] _T_1766;
  wire [15:0] _T_1870;
  wire [15:0] _T_1974;
  wire [15:0] _T_2078;
  wire [15:0] _T_2182;
  wire [15:0] _T_2286;
  wire [15:0] _T_2390;
  wire [15:0] _T_2494;
  wire [15:0] _T_2598;
  wire [15:0] _T_2702;
  wire [15:0] _T_2806;
  wire [15:0] _T_2910;
  wire [15:0] _T_3014;
  wire [15:0] _T_3118;
  wire [15:0] _T_3222;
  wire [15:0] _T_3326;
  wire [15:0] _T_3430;
  wire [15:0] _T_3534;
  wire [15:0] _T_3638;
  wire [15:0] _T_3742;
  wire [15:0] _T_3846;
  wire [15:0] _T_3950;
  wire [15:0] _T_4054;
  wire  _T_4062;
  wire [1:0] _T_4064;
  wire  _T_4065;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_15;
  wire [15:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [15:0] _GEN_20;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_22;
  wire [15:0] _GEN_23;
  wire [15:0] _GEN_24;
  wire [15:0] _GEN_25;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  wire [15:0] _GEN_32;
  wire [15:0] _GEN_33;
  wire [15:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire [15:0] _GEN_36;
  wire [15:0] _GEN_37;
  wire [15:0] _GEN_38;
  wire [15:0] _GEN_39;
  wire [15:0] _GEN_40;
  wire [15:0] _GEN_41;
  wire [15:0] _GEN_42;
  wire [15:0] _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _T_4069;
  wire  _T_4070;
  wire  _T_4072;
  wire [1:0] _T_4075;
  wire  _T_4076;
  wire  _T_4077;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire [1:0] _T_4081;
  wire  _T_4084;
  wire  _T_4086;
  wire [5:0] _T_4090;
  wire [4:0] _T_4091;
  wire  _GEN_49;
  wire [4:0] _GEN_50;
  wire  _GEN_51;
  wire [4:0] _GEN_52;
  wire  _T_4101;
  wire  _T_4106;
  wire  _T_4111;
  wire  _T_4112;
  wire  _T_4114;
  wire [15:0] _GEN_0;
  wire [15:0] _GEN_53;
  wire [15:0] _GEN_54;
  wire [15:0] _GEN_55;
  wire [15:0] _GEN_56;
  wire [15:0] _GEN_57;
  wire [15:0] _GEN_58;
  wire [15:0] _GEN_59;
  wire [15:0] _GEN_60;
  wire [15:0] _GEN_61;
  wire [15:0] _GEN_62;
  wire [15:0] _GEN_63;
  wire [15:0] _GEN_64;
  wire [15:0] _GEN_65;
  wire [15:0] _GEN_66;
  wire [15:0] _GEN_67;
  wire [15:0] _GEN_68;
  wire [15:0] _GEN_69;
  wire [15:0] _GEN_70;
  wire [15:0] _GEN_71;
  wire [15:0] _GEN_72;
  wire [15:0] _GEN_73;
  wire [15:0] _GEN_74;
  wire [15:0] _GEN_75;
  wire [15:0] _GEN_76;
  wire [15:0] _GEN_77;
  wire [15:0] _GEN_78;
  wire [15:0] _GEN_79;
  wire [15:0] _GEN_80;
  wire [15:0] _GEN_81;
  wire [15:0] _GEN_82;
  wire [15:0] _GEN_83;
  wire  _T_4120;
  reg  _T_4123;
  reg [31:0] _RAND_64;
  wire  _T_4125;
  wire [1:0] _T_4127;
  wire  _T_4128;
  wire  _GEN_84;
  reg  _T_4131;
  reg [31:0] _RAND_65;
  wire  _T_4136;
  wire  _T_4137;
  wire  _T_4139;
  wire [1:0] _T_4144;
  wire  _T_4145;
  wire  _T_4146;
  wire [1:0] _T_4150;
  wire  _T_4151;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire  _GEN_90;
  wire  _T_4159;
  wire  _T_4160;
  reg  _T_4163;
  reg [31:0] _RAND_66;
  wire  _T_4165;
  wire [1:0] _T_4167;
  wire  _T_4168;
  wire  _GEN_91;
  reg [15:0] _T_4242_0_0;
  reg [31:0] _RAND_67;
  reg [15:0] _T_4242_0_1;
  reg [31:0] _RAND_68;
  reg [15:0] _T_4242_0_2;
  reg [31:0] _RAND_69;
  reg [15:0] _T_4242_0_3;
  reg [31:0] _RAND_70;
  reg [15:0] _T_4242_0_4;
  reg [31:0] _RAND_71;
  reg [15:0] _T_4242_0_5;
  reg [31:0] _RAND_72;
  reg [15:0] _T_4242_0_6;
  reg [31:0] _RAND_73;
  reg [15:0] _T_4242_0_7;
  reg [31:0] _RAND_74;
  reg [15:0] _T_4242_0_8;
  reg [31:0] _RAND_75;
  reg [15:0] _T_4242_0_9;
  reg [31:0] _RAND_76;
  reg [15:0] _T_4242_0_10;
  reg [31:0] _RAND_77;
  reg [15:0] _T_4242_0_11;
  reg [31:0] _RAND_78;
  reg [15:0] _T_4242_0_12;
  reg [31:0] _RAND_79;
  reg [15:0] _T_4242_0_13;
  reg [31:0] _RAND_80;
  reg [15:0] _T_4242_0_14;
  reg [31:0] _RAND_81;
  reg [15:0] _T_4242_0_15;
  reg [31:0] _RAND_82;
  reg [15:0] _T_4242_0_16;
  reg [31:0] _RAND_83;
  reg [15:0] _T_4242_0_17;
  reg [31:0] _RAND_84;
  reg [15:0] _T_4242_0_18;
  reg [31:0] _RAND_85;
  reg [15:0] _T_4242_0_19;
  reg [31:0] _RAND_86;
  reg [15:0] _T_4242_0_20;
  reg [31:0] _RAND_87;
  reg [15:0] _T_4242_0_21;
  reg [31:0] _RAND_88;
  reg [15:0] _T_4242_0_22;
  reg [31:0] _RAND_89;
  reg [15:0] _T_4242_0_23;
  reg [31:0] _RAND_90;
  reg [15:0] _T_4242_0_24;
  reg [31:0] _RAND_91;
  reg [15:0] _T_4242_0_25;
  reg [31:0] _RAND_92;
  reg [15:0] _T_4242_0_26;
  reg [31:0] _RAND_93;
  reg [15:0] _T_4242_0_27;
  reg [31:0] _RAND_94;
  reg [15:0] _T_4242_0_28;
  reg [31:0] _RAND_95;
  reg [15:0] _T_4242_0_29;
  reg [31:0] _RAND_96;
  reg [15:0] _T_4242_0_30;
  reg [31:0] _RAND_97;
  reg [15:0] _T_4242_0_31;
  reg [31:0] _RAND_98;
  reg [4:0] _T_4461_0;
  reg [31:0] _RAND_99;
  reg  _T_4482_0;
  reg [31:0] _RAND_100;
  reg  _T_4492;
  reg [31:0] _RAND_101;
  wire  _T_4498;
  wire  _T_4499;
  wire  _T_4500;
  wire  _T_4503;
  wire  _T_4504;
  wire [15:0] _T_4608;
  wire [15:0] _T_4712;
  wire [15:0] _T_4816;
  wire [15:0] _T_4920;
  wire [15:0] _T_5024;
  wire [15:0] _T_5128;
  wire [15:0] _T_5232;
  wire [15:0] _T_5336;
  wire [15:0] _T_5440;
  wire [15:0] _T_5544;
  wire [15:0] _T_5648;
  wire [15:0] _T_5752;
  wire [15:0] _T_5856;
  wire [15:0] _T_5960;
  wire [15:0] _T_6064;
  wire [15:0] _T_6168;
  wire [15:0] _T_6272;
  wire [15:0] _T_6376;
  wire [15:0] _T_6480;
  wire [15:0] _T_6584;
  wire [15:0] _T_6688;
  wire [15:0] _T_6792;
  wire [15:0] _T_6896;
  wire [15:0] _T_7000;
  wire [15:0] _T_7104;
  wire [15:0] _T_7208;
  wire [15:0] _T_7312;
  wire [15:0] _T_7416;
  wire [15:0] _T_7520;
  wire [15:0] _T_7624;
  wire [15:0] _T_7728;
  wire [15:0] _T_7832;
  wire  _T_7840;
  wire [1:0] _T_7842;
  wire  _T_7843;
  wire [15:0] _GEN_92;
  wire [15:0] _GEN_93;
  wire [15:0] _GEN_94;
  wire [15:0] _GEN_95;
  wire [15:0] _GEN_96;
  wire [15:0] _GEN_97;
  wire [15:0] _GEN_98;
  wire [15:0] _GEN_99;
  wire [15:0] _GEN_100;
  wire [15:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire [15:0] _GEN_103;
  wire [15:0] _GEN_104;
  wire [15:0] _GEN_105;
  wire [15:0] _GEN_106;
  wire [15:0] _GEN_107;
  wire [15:0] _GEN_108;
  wire [15:0] _GEN_109;
  wire [15:0] _GEN_110;
  wire [15:0] _GEN_111;
  wire [15:0] _GEN_112;
  wire [15:0] _GEN_113;
  wire [15:0] _GEN_114;
  wire [15:0] _GEN_115;
  wire [15:0] _GEN_116;
  wire [15:0] _GEN_117;
  wire [15:0] _GEN_118;
  wire [15:0] _GEN_119;
  wire [15:0] _GEN_120;
  wire [15:0] _GEN_121;
  wire [15:0] _GEN_122;
  wire [15:0] _GEN_123;
  wire  _GEN_124;
  wire  _GEN_125;
  wire  _T_7847;
  wire  _T_7848;
  wire [1:0] _T_7853;
  wire  _T_7854;
  wire  _T_7855;
  wire  _GEN_126;
  wire  _GEN_127;
  wire  _GEN_128;
  wire [1:0] _T_7859;
  wire  _T_7864;
  wire [5:0] _T_7868;
  wire [4:0] _T_7869;
  wire  _GEN_129;
  wire [4:0] _GEN_130;
  wire  _GEN_131;
  wire [4:0] _GEN_132;
  wire  _T_7879;
  wire  _T_7884;
  wire  _T_7889;
  wire  _T_7890;
  wire  _T_7892;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_133;
  wire [15:0] _GEN_134;
  wire [15:0] _GEN_135;
  wire [15:0] _GEN_136;
  wire [15:0] _GEN_137;
  wire [15:0] _GEN_138;
  wire [15:0] _GEN_139;
  wire [15:0] _GEN_140;
  wire [15:0] _GEN_141;
  wire [15:0] _GEN_142;
  wire [15:0] _GEN_143;
  wire [15:0] _GEN_144;
  wire [15:0] _GEN_145;
  wire [15:0] _GEN_146;
  wire [15:0] _GEN_147;
  wire [15:0] _GEN_148;
  wire [15:0] _GEN_149;
  wire [15:0] _GEN_150;
  wire [15:0] _GEN_151;
  wire [15:0] _GEN_152;
  wire [15:0] _GEN_153;
  wire [15:0] _GEN_154;
  wire [15:0] _GEN_155;
  wire [15:0] _GEN_156;
  wire [15:0] _GEN_157;
  wire [15:0] _GEN_158;
  wire [15:0] _GEN_159;
  wire [15:0] _GEN_160;
  wire [15:0] _GEN_161;
  wire [15:0] _GEN_162;
  wire [15:0] _GEN_163;
  wire  _T_7898;
  reg  _T_7901;
  reg [31:0] _RAND_102;
  wire  _T_7903;
  wire [1:0] _T_7905;
  wire  _T_7906;
  wire  _GEN_164;
  reg  _T_7909;
  reg [31:0] _RAND_103;
  reg  _T_7912;
  reg [31:0] _RAND_104;
  reg [15:0] _T_7916_0;
  reg [31:0] _RAND_105;
  reg [15:0] _T_7916_1;
  reg [31:0] _RAND_106;
  reg [15:0] _T_7916_2;
  reg [31:0] _RAND_107;
  reg [15:0] _T_7916_3;
  reg [31:0] _RAND_108;
  reg [15:0] _T_7916_4;
  reg [31:0] _RAND_109;
  reg [15:0] _T_7916_5;
  reg [31:0] _RAND_110;
  reg [15:0] _T_7916_6;
  reg [31:0] _RAND_111;
  reg [15:0] _T_7916_7;
  reg [31:0] _RAND_112;
  reg [15:0] _T_7916_8;
  reg [31:0] _RAND_113;
  reg [15:0] _T_7916_9;
  reg [31:0] _RAND_114;
  reg [15:0] _T_7916_10;
  reg [31:0] _RAND_115;
  reg [15:0] _T_7916_11;
  reg [31:0] _RAND_116;
  reg [15:0] _T_7916_12;
  reg [31:0] _RAND_117;
  reg [15:0] _T_7916_13;
  reg [31:0] _RAND_118;
  reg [15:0] _T_7916_14;
  reg [31:0] _RAND_119;
  reg [15:0] _T_7916_15;
  reg [31:0] _RAND_120;
  reg [15:0] _T_7916_16;
  reg [31:0] _RAND_121;
  reg [15:0] _T_7916_17;
  reg [31:0] _RAND_122;
  reg [15:0] _T_7916_18;
  reg [31:0] _RAND_123;
  reg [15:0] _T_7916_19;
  reg [31:0] _RAND_124;
  reg [15:0] _T_7916_20;
  reg [31:0] _RAND_125;
  reg [15:0] _T_7916_21;
  reg [31:0] _RAND_126;
  reg [15:0] _T_7916_22;
  reg [31:0] _RAND_127;
  reg [15:0] _T_7916_23;
  reg [31:0] _RAND_128;
  reg [15:0] _T_7916_24;
  reg [31:0] _RAND_129;
  reg [15:0] _T_7916_25;
  reg [31:0] _RAND_130;
  reg [15:0] _T_7916_26;
  reg [31:0] _RAND_131;
  reg [15:0] _T_7916_27;
  reg [31:0] _RAND_132;
  reg [15:0] _T_7916_28;
  reg [31:0] _RAND_133;
  reg [15:0] _T_7916_29;
  reg [31:0] _RAND_134;
  reg [15:0] _T_7916_30;
  reg [31:0] _RAND_135;
  reg [15:0] _T_7916_31;
  reg [31:0] _RAND_136;
  reg  _T_7953;
  reg [31:0] _RAND_137;
  wire  _T_7956;
  wire  _T_7958;
  wire  _T_7959;
  wire  _GEN_165;
  wire  _T_7962;
  wire [15:0] _GEN_2;
  wire [15:0] _GEN_166;
  wire [15:0] _GEN_167;
  wire [15:0] _GEN_168;
  wire [15:0] _GEN_169;
  wire [15:0] _GEN_170;
  wire [15:0] _GEN_171;
  wire [15:0] _GEN_172;
  wire [15:0] _GEN_173;
  wire [15:0] _GEN_174;
  wire [15:0] _GEN_175;
  wire [15:0] _GEN_176;
  wire [15:0] _GEN_177;
  wire [15:0] _GEN_178;
  wire [15:0] _GEN_179;
  wire [15:0] _GEN_180;
  wire [15:0] _GEN_181;
  wire [15:0] _GEN_182;
  wire [15:0] _GEN_183;
  wire [15:0] _GEN_184;
  wire [15:0] _GEN_185;
  wire [15:0] _GEN_186;
  wire [15:0] _GEN_187;
  wire [15:0] _GEN_188;
  wire [15:0] _GEN_189;
  wire [15:0] _GEN_190;
  wire [15:0] _GEN_191;
  wire [15:0] _GEN_192;
  wire [15:0] _GEN_193;
  wire [15:0] _GEN_194;
  wire [15:0] _GEN_195;
  wire [15:0] _GEN_196;
  wire [15:0] _GEN_197;
  wire [15:0] _GEN_198;
  wire [15:0] _GEN_199;
  wire [15:0] _GEN_200;
  wire [15:0] _GEN_201;
  wire [15:0] _GEN_202;
  wire [15:0] _GEN_203;
  wire [15:0] _GEN_204;
  wire [15:0] _GEN_205;
  wire [15:0] _GEN_206;
  wire [15:0] _GEN_207;
  wire [15:0] _GEN_208;
  wire [15:0] _GEN_209;
  wire [15:0] _GEN_210;
  wire [15:0] _GEN_211;
  wire [15:0] _GEN_212;
  wire [15:0] _GEN_213;
  wire [15:0] _GEN_214;
  wire [15:0] _GEN_215;
  wire [15:0] _GEN_216;
  wire [15:0] _GEN_217;
  wire [15:0] _GEN_218;
  wire [15:0] _GEN_219;
  wire [15:0] _GEN_220;
  wire [15:0] _GEN_221;
  wire [15:0] _GEN_222;
  wire [15:0] _GEN_223;
  wire [15:0] _GEN_224;
  wire [15:0] _GEN_225;
  wire [15:0] _GEN_226;
  wire [15:0] _GEN_227;
  wire [15:0] _GEN_228;
  wire [15:0] _GEN_229;
  wire  _T_7966;
  wire  _T_7968;
  wire  _T_7969;
  wire  _GEN_230;
  wire  _T_7971;
  wire  _GEN_231;
  wire  _GEN_232;
  wire [31:0] _T_7974;
  wire [31:0] _T_7975;
  wire [63:0] _T_7976;
  wire [31:0] _T_7977;
  wire [31:0] _T_7978;
  wire [63:0] _T_7979;
  wire [127:0] _T_7980;
  wire [31:0] _T_7981;
  wire [31:0] _T_7982;
  wire [63:0] _T_7983;
  wire [31:0] _T_7984;
  wire [31:0] _T_7985;
  wire [63:0] _T_7986;
  wire [127:0] _T_7987;
  wire [255:0] _T_7988;
  wire [31:0] _T_7989;
  wire [31:0] _T_7990;
  wire [63:0] _T_7991;
  wire [31:0] _T_7992;
  wire [31:0] _T_7993;
  wire [63:0] _T_7994;
  wire [127:0] _T_7995;
  wire [31:0] _T_7996;
  wire [31:0] _T_7997;
  wire [63:0] _T_7998;
  wire [31:0] _T_7999;
  wire [31:0] _T_8000;
  wire [63:0] _T_8001;
  wire [127:0] _T_8002;
  wire [255:0] _T_8003;
  wire [511:0] _T_8004;
  wire  _T_8006;
  wire  _T_8008;
  wire  _T_8011;
  wire  _T_8013;
  wire  _T_8014;
  wire  _T_8021;
  wire  _T_8022;
  wire [1:0] _T_8027;
  wire  _T_8028;
  wire  _T_8029;
  wire  _GEN_233;
  wire  _GEN_234;
  wire  _GEN_235;
  wire  _GEN_236;
  reg  _T_8035;
  reg [31:0] _RAND_138;
  wire  _T_8037;
  wire [1:0] _T_8039;
  wire  _T_8040;
  wire  _GEN_237;
  reg  _T_8043;
  reg [31:0] _RAND_139;
  reg  _T_8046;
  reg [31:0] _RAND_140;
  reg [15:0] _T_8050_0;
  reg [31:0] _RAND_141;
  reg [15:0] _T_8050_1;
  reg [31:0] _RAND_142;
  reg [15:0] _T_8050_2;
  reg [31:0] _RAND_143;
  reg [15:0] _T_8050_3;
  reg [31:0] _RAND_144;
  reg [15:0] _T_8050_4;
  reg [31:0] _RAND_145;
  reg [15:0] _T_8050_5;
  reg [31:0] _RAND_146;
  reg [15:0] _T_8050_6;
  reg [31:0] _RAND_147;
  reg [15:0] _T_8050_7;
  reg [31:0] _RAND_148;
  reg [15:0] _T_8050_8;
  reg [31:0] _RAND_149;
  reg [15:0] _T_8050_9;
  reg [31:0] _RAND_150;
  reg [15:0] _T_8050_10;
  reg [31:0] _RAND_151;
  reg [15:0] _T_8050_11;
  reg [31:0] _RAND_152;
  reg [15:0] _T_8050_12;
  reg [31:0] _RAND_153;
  reg [15:0] _T_8050_13;
  reg [31:0] _RAND_154;
  reg [15:0] _T_8050_14;
  reg [31:0] _RAND_155;
  reg [15:0] _T_8050_15;
  reg [31:0] _RAND_156;
  reg [15:0] _T_8050_16;
  reg [31:0] _RAND_157;
  reg [15:0] _T_8050_17;
  reg [31:0] _RAND_158;
  reg [15:0] _T_8050_18;
  reg [31:0] _RAND_159;
  reg [15:0] _T_8050_19;
  reg [31:0] _RAND_160;
  reg [15:0] _T_8050_20;
  reg [31:0] _RAND_161;
  reg [15:0] _T_8050_21;
  reg [31:0] _RAND_162;
  reg [15:0] _T_8050_22;
  reg [31:0] _RAND_163;
  reg [15:0] _T_8050_23;
  reg [31:0] _RAND_164;
  reg [15:0] _T_8050_24;
  reg [31:0] _RAND_165;
  reg [15:0] _T_8050_25;
  reg [31:0] _RAND_166;
  reg [15:0] _T_8050_26;
  reg [31:0] _RAND_167;
  reg [15:0] _T_8050_27;
  reg [31:0] _RAND_168;
  reg [15:0] _T_8050_28;
  reg [31:0] _RAND_169;
  reg [15:0] _T_8050_29;
  reg [31:0] _RAND_170;
  reg [15:0] _T_8050_30;
  reg [31:0] _RAND_171;
  reg [15:0] _T_8050_31;
  reg [31:0] _RAND_172;
  reg  _T_8087;
  reg [31:0] _RAND_173;
  wire  _T_8090;
  wire  _T_8092;
  wire  _T_8093;
  wire  _GEN_238;
  wire  _T_8096;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_239;
  wire [15:0] _GEN_240;
  wire [15:0] _GEN_241;
  wire [15:0] _GEN_242;
  wire [15:0] _GEN_243;
  wire [15:0] _GEN_244;
  wire [15:0] _GEN_245;
  wire [15:0] _GEN_246;
  wire [15:0] _GEN_247;
  wire [15:0] _GEN_248;
  wire [15:0] _GEN_249;
  wire [15:0] _GEN_250;
  wire [15:0] _GEN_251;
  wire [15:0] _GEN_252;
  wire [15:0] _GEN_253;
  wire [15:0] _GEN_254;
  wire [15:0] _GEN_255;
  wire [15:0] _GEN_256;
  wire [15:0] _GEN_257;
  wire [15:0] _GEN_258;
  wire [15:0] _GEN_259;
  wire [15:0] _GEN_260;
  wire [15:0] _GEN_261;
  wire [15:0] _GEN_262;
  wire [15:0] _GEN_263;
  wire [15:0] _GEN_264;
  wire [15:0] _GEN_265;
  wire [15:0] _GEN_266;
  wire [15:0] _GEN_267;
  wire [15:0] _GEN_268;
  wire [15:0] _GEN_269;
  wire [15:0] _GEN_270;
  wire [15:0] _GEN_271;
  wire [15:0] _GEN_272;
  wire [15:0] _GEN_273;
  wire [15:0] _GEN_274;
  wire [15:0] _GEN_275;
  wire [15:0] _GEN_276;
  wire [15:0] _GEN_277;
  wire [15:0] _GEN_278;
  wire [15:0] _GEN_279;
  wire [15:0] _GEN_280;
  wire [15:0] _GEN_281;
  wire [15:0] _GEN_282;
  wire [15:0] _GEN_283;
  wire [15:0] _GEN_284;
  wire [15:0] _GEN_285;
  wire [15:0] _GEN_286;
  wire [15:0] _GEN_287;
  wire [15:0] _GEN_288;
  wire [15:0] _GEN_289;
  wire [15:0] _GEN_290;
  wire [15:0] _GEN_291;
  wire [15:0] _GEN_292;
  wire [15:0] _GEN_293;
  wire [15:0] _GEN_294;
  wire [15:0] _GEN_295;
  wire [15:0] _GEN_296;
  wire [15:0] _GEN_297;
  wire [15:0] _GEN_298;
  wire [15:0] _GEN_299;
  wire [15:0] _GEN_300;
  wire [15:0] _GEN_301;
  wire [15:0] _GEN_302;
  wire  _T_8100;
  wire  _T_8102;
  wire  _T_8103;
  wire  _GEN_303;
  wire  _T_8105;
  wire  _GEN_304;
  wire  _GEN_305;
  wire [31:0] _T_8108;
  wire [31:0] _T_8109;
  wire [63:0] _T_8110;
  wire [31:0] _T_8111;
  wire [31:0] _T_8112;
  wire [63:0] _T_8113;
  wire [127:0] _T_8114;
  wire [31:0] _T_8115;
  wire [31:0] _T_8116;
  wire [63:0] _T_8117;
  wire [31:0] _T_8118;
  wire [31:0] _T_8119;
  wire [63:0] _T_8120;
  wire [127:0] _T_8121;
  wire [255:0] _T_8122;
  wire [31:0] _T_8123;
  wire [31:0] _T_8124;
  wire [63:0] _T_8125;
  wire [31:0] _T_8126;
  wire [31:0] _T_8127;
  wire [63:0] _T_8128;
  wire [127:0] _T_8129;
  wire [31:0] _T_8130;
  wire [31:0] _T_8131;
  wire [63:0] _T_8132;
  wire [31:0] _T_8133;
  wire [31:0] _T_8134;
  wire [63:0] _T_8135;
  wire [127:0] _T_8136;
  wire [255:0] _T_8137;
  wire [511:0] _T_8138;
  wire  _T_8142;
  wire  _T_8145;
  wire  _T_8147;
  wire  _T_8148;
  wire  _T_8155;
  wire  _T_8156;
  wire [1:0] _T_8161;
  wire  _T_8162;
  wire  _T_8163;
  wire  _GEN_306;
  wire  _GEN_307;
  wire  _GEN_308;
  wire  _GEN_309;
  wire  cumFinished;
  StreamingCore StreamingCore (
    .clock(StreamingCore_clock),
    .reset(StreamingCore_reset),
    .io_inputMemAddr(StreamingCore_io_inputMemAddr),
    .io_inputMemAddrConsumed(StreamingCore_io_inputMemAddrConsumed),
    .io_inputMemBlock(StreamingCore_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_io_outputMemBlockReady),
    .io_inputAddrsIgnore(StreamingCore_io_inputAddrsIgnore),
    .io_inputBlocksFinished(StreamingCore_io_inputBlocksFinished),
    .io_outputFinished(StreamingCore_io_outputFinished)
  );
  StreamingCore_1 StreamingCore_1 (
    .clock(StreamingCore_1_clock),
    .reset(StreamingCore_1_reset),
    .io_inputMemAddr(StreamingCore_1_io_inputMemAddr),
    .io_inputMemAddrConsumed(StreamingCore_1_io_inputMemAddrConsumed),
    .io_inputMemBlock(StreamingCore_1_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_1_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_1_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_1_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_1_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_1_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_1_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_1_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_1_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_1_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_1_io_outputMemBlockReady),
    .io_inputAddrsIgnore(StreamingCore_1_io_inputAddrsIgnore),
    .io_inputBlocksFinished(StreamingCore_1_io_inputBlocksFinished),
    .io_outputFinished(StreamingCore_1_io_outputFinished)
  );
  assign _T_347 = _T_345 != 1'h1;
  assign _T_349 = _T_345 + 1'h1;
  assign _T_350 = _T_349[0:0];
  assign _GEN_4 = _T_347 ? _T_350 : _T_345;
  assign _T_358 = io_inputMemAddrReadys_0 | _T_277_0;
  assign _T_359 = _T_345 & _T_358;
  assign _T_361 = _T_353 == 1'h0;
  assign _T_363 = _T_239 == 1'h0;
  assign _T_366 = _T_239 + 1'h1;
  assign _T_367 = _T_366[0:0];
  assign _T_368 = _T_363 ? 1'h0 : _T_367;
  assign _T_372 = _T_353 + 1'h1;
  assign _T_373 = _T_372[0:0];
  assign _GEN_5 = _T_361 ? _T_368 : _T_239;
  assign _GEN_6 = _T_361 ? 1'h0 : _GEN_4;
  assign _GEN_7 = _T_361 ? 1'h0 : _T_373;
  assign _GEN_8 = _T_359 ? _GEN_5 : _T_239;
  assign _GEN_9 = _T_359 ? _GEN_6 : _GEN_4;
  assign _GEN_10 = _T_359 ? _GEN_7 : _T_353;
  assign _T_381 = _T_277_0 == 1'h0;
  assign _T_382 = _T_345 & _T_381;
  assign _T_387 = _T_385 != 1'h1;
  assign _T_389 = _T_385 + 1'h1;
  assign _T_390 = _T_389[0:0];
  assign _GEN_11 = _T_387 ? _T_390 : _T_385;
  assign _T_720 = _T_714 == 1'h0;
  assign _T_721 = _T_385 & _T_720;
  assign _T_722 = io_inputMemBlockReadys_0 & io_inputMemBlockValids_0;
  assign _T_725 = _T_722 | _T_283_0;
  assign _T_726 = _T_721 & _T_725;
  assign _T_830 = io_inputMemBlocks_0[15:0];
  assign _T_934 = io_inputMemBlocks_0[31:16];
  assign _T_1038 = io_inputMemBlocks_0[47:32];
  assign _T_1142 = io_inputMemBlocks_0[63:48];
  assign _T_1246 = io_inputMemBlocks_0[79:64];
  assign _T_1350 = io_inputMemBlocks_0[95:80];
  assign _T_1454 = io_inputMemBlocks_0[111:96];
  assign _T_1558 = io_inputMemBlocks_0[127:112];
  assign _T_1662 = io_inputMemBlocks_0[143:128];
  assign _T_1766 = io_inputMemBlocks_0[159:144];
  assign _T_1870 = io_inputMemBlocks_0[175:160];
  assign _T_1974 = io_inputMemBlocks_0[191:176];
  assign _T_2078 = io_inputMemBlocks_0[207:192];
  assign _T_2182 = io_inputMemBlocks_0[223:208];
  assign _T_2286 = io_inputMemBlocks_0[239:224];
  assign _T_2390 = io_inputMemBlocks_0[255:240];
  assign _T_2494 = io_inputMemBlocks_0[271:256];
  assign _T_2598 = io_inputMemBlocks_0[287:272];
  assign _T_2702 = io_inputMemBlocks_0[303:288];
  assign _T_2806 = io_inputMemBlocks_0[319:304];
  assign _T_2910 = io_inputMemBlocks_0[335:320];
  assign _T_3014 = io_inputMemBlocks_0[351:336];
  assign _T_3118 = io_inputMemBlocks_0[367:352];
  assign _T_3222 = io_inputMemBlocks_0[383:368];
  assign _T_3326 = io_inputMemBlocks_0[399:384];
  assign _T_3430 = io_inputMemBlocks_0[415:400];
  assign _T_3534 = io_inputMemBlocks_0[431:416];
  assign _T_3638 = io_inputMemBlocks_0[447:432];
  assign _T_3742 = io_inputMemBlocks_0[463:448];
  assign _T_3846 = io_inputMemBlocks_0[479:464];
  assign _T_3950 = io_inputMemBlocks_0[495:480];
  assign _T_4054 = io_inputMemBlocks_0[511:496];
  assign _T_4062 = _T_283_0 == 1'h0;
  assign _T_4064 = _T_714 + 1'h1;
  assign _T_4065 = _T_4064[0:0];
  assign _GEN_12 = _T_726 ? _T_830 : _T_464_0_0;
  assign _GEN_13 = _T_726 ? _T_934 : _T_464_0_1;
  assign _GEN_14 = _T_726 ? _T_1038 : _T_464_0_2;
  assign _GEN_15 = _T_726 ? _T_1142 : _T_464_0_3;
  assign _GEN_16 = _T_726 ? _T_1246 : _T_464_0_4;
  assign _GEN_17 = _T_726 ? _T_1350 : _T_464_0_5;
  assign _GEN_18 = _T_726 ? _T_1454 : _T_464_0_6;
  assign _GEN_19 = _T_726 ? _T_1558 : _T_464_0_7;
  assign _GEN_20 = _T_726 ? _T_1662 : _T_464_0_8;
  assign _GEN_21 = _T_726 ? _T_1766 : _T_464_0_9;
  assign _GEN_22 = _T_726 ? _T_1870 : _T_464_0_10;
  assign _GEN_23 = _T_726 ? _T_1974 : _T_464_0_11;
  assign _GEN_24 = _T_726 ? _T_2078 : _T_464_0_12;
  assign _GEN_25 = _T_726 ? _T_2182 : _T_464_0_13;
  assign _GEN_26 = _T_726 ? _T_2286 : _T_464_0_14;
  assign _GEN_27 = _T_726 ? _T_2390 : _T_464_0_15;
  assign _GEN_28 = _T_726 ? _T_2494 : _T_464_0_16;
  assign _GEN_29 = _T_726 ? _T_2598 : _T_464_0_17;
  assign _GEN_30 = _T_726 ? _T_2702 : _T_464_0_18;
  assign _GEN_31 = _T_726 ? _T_2806 : _T_464_0_19;
  assign _GEN_32 = _T_726 ? _T_2910 : _T_464_0_20;
  assign _GEN_33 = _T_726 ? _T_3014 : _T_464_0_21;
  assign _GEN_34 = _T_726 ? _T_3118 : _T_464_0_22;
  assign _GEN_35 = _T_726 ? _T_3222 : _T_464_0_23;
  assign _GEN_36 = _T_726 ? _T_3326 : _T_464_0_24;
  assign _GEN_37 = _T_726 ? _T_3430 : _T_464_0_25;
  assign _GEN_38 = _T_726 ? _T_3534 : _T_464_0_26;
  assign _GEN_39 = _T_726 ? _T_3638 : _T_464_0_27;
  assign _GEN_40 = _T_726 ? _T_3742 : _T_464_0_28;
  assign _GEN_41 = _T_726 ? _T_3846 : _T_464_0_29;
  assign _GEN_42 = _T_726 ? _T_3950 : _T_464_0_30;
  assign _GEN_43 = _T_726 ? _T_4054 : _T_464_0_31;
  assign _GEN_44 = _T_726 ? _T_4062 : _T_704_0;
  assign _GEN_45 = _T_726 ? _T_4065 : _T_714;
  assign _T_4069 = _T_704_0 == 1'h0;
  assign _T_4070 = _T_714 & _T_4069;
  assign _T_4072 = _T_242 == 1'h0;
  assign _T_4075 = _T_242 + 1'h1;
  assign _T_4076 = _T_4075[0:0];
  assign _T_4077 = _T_4072 ? 1'h0 : _T_4076;
  assign _GEN_46 = _T_4070 ? _T_4077 : _T_242;
  assign _GEN_47 = _T_4070 ? 1'h0 : _GEN_11;
  assign _GEN_48 = _T_4070 ? 1'h0 : _GEN_45;
  assign _T_4081 = {_T_242,_T_714};
  assign _T_4084 = reset == 1'h0;
  assign _T_4086 = _T_683_0 == 5'h1f;
  assign _T_4090 = _T_683_0 + 5'h1;
  assign _T_4091 = _T_4090[4:0];
  assign _GEN_49 = _T_4086 ? 1'h0 : _GEN_44;
  assign _GEN_50 = _T_4086 ? 5'h0 : _T_4091;
  assign _GEN_51 = _T_704_0 ? _GEN_49 : _GEN_44;
  assign _GEN_52 = _T_704_0 ? _GEN_50 : _T_683_0;
  assign _T_4101 = _T_721 & _T_271_0;
  assign _T_4106 = _T_4101 & _T_4062;
  assign _T_4111 = _T_361 & io_inputMemAddrReadys_0;
  assign _T_4112 = _T_4111 & io_inputMemAddrValids_0;
  assign _T_4114 = _T_363 ? _T_4112 : 1'h0;
  assign _GEN_53 = 5'h1 == _T_683_0 ? _T_464_0_1 : _T_464_0_0;
  assign _GEN_54 = 5'h2 == _T_683_0 ? _T_464_0_2 : _GEN_53;
  assign _GEN_55 = 5'h3 == _T_683_0 ? _T_464_0_3 : _GEN_54;
  assign _GEN_56 = 5'h4 == _T_683_0 ? _T_464_0_4 : _GEN_55;
  assign _GEN_57 = 5'h5 == _T_683_0 ? _T_464_0_5 : _GEN_56;
  assign _GEN_58 = 5'h6 == _T_683_0 ? _T_464_0_6 : _GEN_57;
  assign _GEN_59 = 5'h7 == _T_683_0 ? _T_464_0_7 : _GEN_58;
  assign _GEN_60 = 5'h8 == _T_683_0 ? _T_464_0_8 : _GEN_59;
  assign _GEN_61 = 5'h9 == _T_683_0 ? _T_464_0_9 : _GEN_60;
  assign _GEN_62 = 5'ha == _T_683_0 ? _T_464_0_10 : _GEN_61;
  assign _GEN_63 = 5'hb == _T_683_0 ? _T_464_0_11 : _GEN_62;
  assign _GEN_64 = 5'hc == _T_683_0 ? _T_464_0_12 : _GEN_63;
  assign _GEN_65 = 5'hd == _T_683_0 ? _T_464_0_13 : _GEN_64;
  assign _GEN_66 = 5'he == _T_683_0 ? _T_464_0_14 : _GEN_65;
  assign _GEN_67 = 5'hf == _T_683_0 ? _T_464_0_15 : _GEN_66;
  assign _GEN_68 = 5'h10 == _T_683_0 ? _T_464_0_16 : _GEN_67;
  assign _GEN_69 = 5'h11 == _T_683_0 ? _T_464_0_17 : _GEN_68;
  assign _GEN_70 = 5'h12 == _T_683_0 ? _T_464_0_18 : _GEN_69;
  assign _GEN_71 = 5'h13 == _T_683_0 ? _T_464_0_19 : _GEN_70;
  assign _GEN_72 = 5'h14 == _T_683_0 ? _T_464_0_20 : _GEN_71;
  assign _GEN_73 = 5'h15 == _T_683_0 ? _T_464_0_21 : _GEN_72;
  assign _GEN_74 = 5'h16 == _T_683_0 ? _T_464_0_22 : _GEN_73;
  assign _GEN_75 = 5'h17 == _T_683_0 ? _T_464_0_23 : _GEN_74;
  assign _GEN_76 = 5'h18 == _T_683_0 ? _T_464_0_24 : _GEN_75;
  assign _GEN_77 = 5'h19 == _T_683_0 ? _T_464_0_25 : _GEN_76;
  assign _GEN_78 = 5'h1a == _T_683_0 ? _T_464_0_26 : _GEN_77;
  assign _GEN_79 = 5'h1b == _T_683_0 ? _T_464_0_27 : _GEN_78;
  assign _GEN_80 = 5'h1c == _T_683_0 ? _T_464_0_28 : _GEN_79;
  assign _GEN_81 = 5'h1d == _T_683_0 ? _T_464_0_29 : _GEN_80;
  assign _GEN_82 = 5'h1e == _T_683_0 ? _T_464_0_30 : _GEN_81;
  assign _GEN_83 = 5'h1f == _T_683_0 ? _T_464_0_31 : _GEN_82;
  assign _T_4120 = _T_4072 ? _T_704_0 : 1'h0;
  assign _T_4125 = _T_4123 != 1'h1;
  assign _T_4127 = _T_4123 + 1'h1;
  assign _T_4128 = _T_4127[0:0];
  assign _GEN_84 = _T_4125 ? _T_4128 : _T_4123;
  assign _T_4136 = io_inputMemAddrReadys_1 | _T_309_0;
  assign _T_4137 = _T_4123 & _T_4136;
  assign _T_4139 = _T_4131 == 1'h0;
  assign _T_4144 = _T_245 + 1'h1;
  assign _T_4145 = _T_4144[0:0];
  assign _T_4146 = _T_245 ? 1'h1 : _T_4145;
  assign _T_4150 = _T_4131 + 1'h1;
  assign _T_4151 = _T_4150[0:0];
  assign _GEN_85 = _T_4139 ? _T_4146 : _T_245;
  assign _GEN_86 = _T_4139 ? 1'h0 : _GEN_84;
  assign _GEN_87 = _T_4139 ? 1'h0 : _T_4151;
  assign _GEN_88 = _T_4137 ? _GEN_85 : _T_245;
  assign _GEN_89 = _T_4137 ? _GEN_86 : _GEN_84;
  assign _GEN_90 = _T_4137 ? _GEN_87 : _T_4131;
  assign _T_4159 = _T_309_0 == 1'h0;
  assign _T_4160 = _T_4123 & _T_4159;
  assign _T_4165 = _T_4163 != 1'h1;
  assign _T_4167 = _T_4163 + 1'h1;
  assign _T_4168 = _T_4167[0:0];
  assign _GEN_91 = _T_4165 ? _T_4168 : _T_4163;
  assign _T_4498 = _T_4492 == 1'h0;
  assign _T_4499 = _T_4163 & _T_4498;
  assign _T_4500 = io_inputMemBlockReadys_1 & io_inputMemBlockValids_1;
  assign _T_4503 = _T_4500 | _T_315_0;
  assign _T_4504 = _T_4499 & _T_4503;
  assign _T_4608 = io_inputMemBlocks_1[15:0];
  assign _T_4712 = io_inputMemBlocks_1[31:16];
  assign _T_4816 = io_inputMemBlocks_1[47:32];
  assign _T_4920 = io_inputMemBlocks_1[63:48];
  assign _T_5024 = io_inputMemBlocks_1[79:64];
  assign _T_5128 = io_inputMemBlocks_1[95:80];
  assign _T_5232 = io_inputMemBlocks_1[111:96];
  assign _T_5336 = io_inputMemBlocks_1[127:112];
  assign _T_5440 = io_inputMemBlocks_1[143:128];
  assign _T_5544 = io_inputMemBlocks_1[159:144];
  assign _T_5648 = io_inputMemBlocks_1[175:160];
  assign _T_5752 = io_inputMemBlocks_1[191:176];
  assign _T_5856 = io_inputMemBlocks_1[207:192];
  assign _T_5960 = io_inputMemBlocks_1[223:208];
  assign _T_6064 = io_inputMemBlocks_1[239:224];
  assign _T_6168 = io_inputMemBlocks_1[255:240];
  assign _T_6272 = io_inputMemBlocks_1[271:256];
  assign _T_6376 = io_inputMemBlocks_1[287:272];
  assign _T_6480 = io_inputMemBlocks_1[303:288];
  assign _T_6584 = io_inputMemBlocks_1[319:304];
  assign _T_6688 = io_inputMemBlocks_1[335:320];
  assign _T_6792 = io_inputMemBlocks_1[351:336];
  assign _T_6896 = io_inputMemBlocks_1[367:352];
  assign _T_7000 = io_inputMemBlocks_1[383:368];
  assign _T_7104 = io_inputMemBlocks_1[399:384];
  assign _T_7208 = io_inputMemBlocks_1[415:400];
  assign _T_7312 = io_inputMemBlocks_1[431:416];
  assign _T_7416 = io_inputMemBlocks_1[447:432];
  assign _T_7520 = io_inputMemBlocks_1[463:448];
  assign _T_7624 = io_inputMemBlocks_1[479:464];
  assign _T_7728 = io_inputMemBlocks_1[495:480];
  assign _T_7832 = io_inputMemBlocks_1[511:496];
  assign _T_7840 = _T_315_0 == 1'h0;
  assign _T_7842 = _T_4492 + 1'h1;
  assign _T_7843 = _T_7842[0:0];
  assign _GEN_92 = _T_4504 ? _T_4608 : _T_4242_0_0;
  assign _GEN_93 = _T_4504 ? _T_4712 : _T_4242_0_1;
  assign _GEN_94 = _T_4504 ? _T_4816 : _T_4242_0_2;
  assign _GEN_95 = _T_4504 ? _T_4920 : _T_4242_0_3;
  assign _GEN_96 = _T_4504 ? _T_5024 : _T_4242_0_4;
  assign _GEN_97 = _T_4504 ? _T_5128 : _T_4242_0_5;
  assign _GEN_98 = _T_4504 ? _T_5232 : _T_4242_0_6;
  assign _GEN_99 = _T_4504 ? _T_5336 : _T_4242_0_7;
  assign _GEN_100 = _T_4504 ? _T_5440 : _T_4242_0_8;
  assign _GEN_101 = _T_4504 ? _T_5544 : _T_4242_0_9;
  assign _GEN_102 = _T_4504 ? _T_5648 : _T_4242_0_10;
  assign _GEN_103 = _T_4504 ? _T_5752 : _T_4242_0_11;
  assign _GEN_104 = _T_4504 ? _T_5856 : _T_4242_0_12;
  assign _GEN_105 = _T_4504 ? _T_5960 : _T_4242_0_13;
  assign _GEN_106 = _T_4504 ? _T_6064 : _T_4242_0_14;
  assign _GEN_107 = _T_4504 ? _T_6168 : _T_4242_0_15;
  assign _GEN_108 = _T_4504 ? _T_6272 : _T_4242_0_16;
  assign _GEN_109 = _T_4504 ? _T_6376 : _T_4242_0_17;
  assign _GEN_110 = _T_4504 ? _T_6480 : _T_4242_0_18;
  assign _GEN_111 = _T_4504 ? _T_6584 : _T_4242_0_19;
  assign _GEN_112 = _T_4504 ? _T_6688 : _T_4242_0_20;
  assign _GEN_113 = _T_4504 ? _T_6792 : _T_4242_0_21;
  assign _GEN_114 = _T_4504 ? _T_6896 : _T_4242_0_22;
  assign _GEN_115 = _T_4504 ? _T_7000 : _T_4242_0_23;
  assign _GEN_116 = _T_4504 ? _T_7104 : _T_4242_0_24;
  assign _GEN_117 = _T_4504 ? _T_7208 : _T_4242_0_25;
  assign _GEN_118 = _T_4504 ? _T_7312 : _T_4242_0_26;
  assign _GEN_119 = _T_4504 ? _T_7416 : _T_4242_0_27;
  assign _GEN_120 = _T_4504 ? _T_7520 : _T_4242_0_28;
  assign _GEN_121 = _T_4504 ? _T_7624 : _T_4242_0_29;
  assign _GEN_122 = _T_4504 ? _T_7728 : _T_4242_0_30;
  assign _GEN_123 = _T_4504 ? _T_7832 : _T_4242_0_31;
  assign _GEN_124 = _T_4504 ? _T_7840 : _T_4482_0;
  assign _GEN_125 = _T_4504 ? _T_7843 : _T_4492;
  assign _T_7847 = _T_4482_0 == 1'h0;
  assign _T_7848 = _T_4492 & _T_7847;
  assign _T_7853 = _T_248 + 1'h1;
  assign _T_7854 = _T_7853[0:0];
  assign _T_7855 = _T_248 ? 1'h1 : _T_7854;
  assign _GEN_126 = _T_7848 ? _T_7855 : _T_248;
  assign _GEN_127 = _T_7848 ? 1'h0 : _GEN_91;
  assign _GEN_128 = _T_7848 ? 1'h0 : _GEN_125;
  assign _T_7859 = {_T_248,_T_4492};
  assign _T_7864 = _T_4461_0 == 5'h1f;
  assign _T_7868 = _T_4461_0 + 5'h1;
  assign _T_7869 = _T_7868[4:0];
  assign _GEN_129 = _T_7864 ? 1'h0 : _GEN_124;
  assign _GEN_130 = _T_7864 ? 5'h0 : _T_7869;
  assign _GEN_131 = _T_4482_0 ? _GEN_129 : _GEN_124;
  assign _GEN_132 = _T_4482_0 ? _GEN_130 : _T_4461_0;
  assign _T_7879 = _T_4499 & _T_303_0;
  assign _T_7884 = _T_7879 & _T_7840;
  assign _T_7889 = _T_4139 & io_inputMemAddrReadys_1;
  assign _T_7890 = _T_7889 & io_inputMemAddrValids_1;
  assign _T_7892 = _T_245 ? _T_7890 : 1'h0;
  assign _GEN_133 = 5'h1 == _T_4461_0 ? _T_4242_0_1 : _T_4242_0_0;
  assign _GEN_134 = 5'h2 == _T_4461_0 ? _T_4242_0_2 : _GEN_133;
  assign _GEN_135 = 5'h3 == _T_4461_0 ? _T_4242_0_3 : _GEN_134;
  assign _GEN_136 = 5'h4 == _T_4461_0 ? _T_4242_0_4 : _GEN_135;
  assign _GEN_137 = 5'h5 == _T_4461_0 ? _T_4242_0_5 : _GEN_136;
  assign _GEN_138 = 5'h6 == _T_4461_0 ? _T_4242_0_6 : _GEN_137;
  assign _GEN_139 = 5'h7 == _T_4461_0 ? _T_4242_0_7 : _GEN_138;
  assign _GEN_140 = 5'h8 == _T_4461_0 ? _T_4242_0_8 : _GEN_139;
  assign _GEN_141 = 5'h9 == _T_4461_0 ? _T_4242_0_9 : _GEN_140;
  assign _GEN_142 = 5'ha == _T_4461_0 ? _T_4242_0_10 : _GEN_141;
  assign _GEN_143 = 5'hb == _T_4461_0 ? _T_4242_0_11 : _GEN_142;
  assign _GEN_144 = 5'hc == _T_4461_0 ? _T_4242_0_12 : _GEN_143;
  assign _GEN_145 = 5'hd == _T_4461_0 ? _T_4242_0_13 : _GEN_144;
  assign _GEN_146 = 5'he == _T_4461_0 ? _T_4242_0_14 : _GEN_145;
  assign _GEN_147 = 5'hf == _T_4461_0 ? _T_4242_0_15 : _GEN_146;
  assign _GEN_148 = 5'h10 == _T_4461_0 ? _T_4242_0_16 : _GEN_147;
  assign _GEN_149 = 5'h11 == _T_4461_0 ? _T_4242_0_17 : _GEN_148;
  assign _GEN_150 = 5'h12 == _T_4461_0 ? _T_4242_0_18 : _GEN_149;
  assign _GEN_151 = 5'h13 == _T_4461_0 ? _T_4242_0_19 : _GEN_150;
  assign _GEN_152 = 5'h14 == _T_4461_0 ? _T_4242_0_20 : _GEN_151;
  assign _GEN_153 = 5'h15 == _T_4461_0 ? _T_4242_0_21 : _GEN_152;
  assign _GEN_154 = 5'h16 == _T_4461_0 ? _T_4242_0_22 : _GEN_153;
  assign _GEN_155 = 5'h17 == _T_4461_0 ? _T_4242_0_23 : _GEN_154;
  assign _GEN_156 = 5'h18 == _T_4461_0 ? _T_4242_0_24 : _GEN_155;
  assign _GEN_157 = 5'h19 == _T_4461_0 ? _T_4242_0_25 : _GEN_156;
  assign _GEN_158 = 5'h1a == _T_4461_0 ? _T_4242_0_26 : _GEN_157;
  assign _GEN_159 = 5'h1b == _T_4461_0 ? _T_4242_0_27 : _GEN_158;
  assign _GEN_160 = 5'h1c == _T_4461_0 ? _T_4242_0_28 : _GEN_159;
  assign _GEN_161 = 5'h1d == _T_4461_0 ? _T_4242_0_29 : _GEN_160;
  assign _GEN_162 = 5'h1e == _T_4461_0 ? _T_4242_0_30 : _GEN_161;
  assign _GEN_163 = 5'h1f == _T_4461_0 ? _T_4242_0_31 : _GEN_162;
  assign _T_7898 = _T_248 ? _T_4482_0 : 1'h0;
  assign _T_7903 = _T_7901 != 1'h1;
  assign _T_7905 = _T_7901 + 1'h1;
  assign _T_7906 = _T_7905[0:0];
  assign _GEN_164 = _T_7903 ? _T_7906 : _T_7901;
  assign _T_7956 = _T_7901 & _T_324;
  assign _T_7958 = _T_328 == 5'h1f;
  assign _T_7959 = _T_7956 & _T_7958;
  assign _GEN_165 = _T_7959 ? 1'h1 : _T_7953;
  assign _T_7962 = _T_7953 == 1'h0;
  assign _GEN_166 = 5'h0 == _T_328 ? _GEN_2 : _T_7916_0;
  assign _GEN_167 = 5'h1 == _T_328 ? _GEN_2 : _T_7916_1;
  assign _GEN_168 = 5'h2 == _T_328 ? _GEN_2 : _T_7916_2;
  assign _GEN_169 = 5'h3 == _T_328 ? _GEN_2 : _T_7916_3;
  assign _GEN_170 = 5'h4 == _T_328 ? _GEN_2 : _T_7916_4;
  assign _GEN_171 = 5'h5 == _T_328 ? _GEN_2 : _T_7916_5;
  assign _GEN_172 = 5'h6 == _T_328 ? _GEN_2 : _T_7916_6;
  assign _GEN_173 = 5'h7 == _T_328 ? _GEN_2 : _T_7916_7;
  assign _GEN_174 = 5'h8 == _T_328 ? _GEN_2 : _T_7916_8;
  assign _GEN_175 = 5'h9 == _T_328 ? _GEN_2 : _T_7916_9;
  assign _GEN_176 = 5'ha == _T_328 ? _GEN_2 : _T_7916_10;
  assign _GEN_177 = 5'hb == _T_328 ? _GEN_2 : _T_7916_11;
  assign _GEN_178 = 5'hc == _T_328 ? _GEN_2 : _T_7916_12;
  assign _GEN_179 = 5'hd == _T_328 ? _GEN_2 : _T_7916_13;
  assign _GEN_180 = 5'he == _T_328 ? _GEN_2 : _T_7916_14;
  assign _GEN_181 = 5'hf == _T_328 ? _GEN_2 : _T_7916_15;
  assign _GEN_182 = 5'h10 == _T_328 ? _GEN_2 : _T_7916_16;
  assign _GEN_183 = 5'h11 == _T_328 ? _GEN_2 : _T_7916_17;
  assign _GEN_184 = 5'h12 == _T_328 ? _GEN_2 : _T_7916_18;
  assign _GEN_185 = 5'h13 == _T_328 ? _GEN_2 : _T_7916_19;
  assign _GEN_186 = 5'h14 == _T_328 ? _GEN_2 : _T_7916_20;
  assign _GEN_187 = 5'h15 == _T_328 ? _GEN_2 : _T_7916_21;
  assign _GEN_188 = 5'h16 == _T_328 ? _GEN_2 : _T_7916_22;
  assign _GEN_189 = 5'h17 == _T_328 ? _GEN_2 : _T_7916_23;
  assign _GEN_190 = 5'h18 == _T_328 ? _GEN_2 : _T_7916_24;
  assign _GEN_191 = 5'h19 == _T_328 ? _GEN_2 : _T_7916_25;
  assign _GEN_192 = 5'h1a == _T_328 ? _GEN_2 : _T_7916_26;
  assign _GEN_193 = 5'h1b == _T_328 ? _GEN_2 : _T_7916_27;
  assign _GEN_194 = 5'h1c == _T_328 ? _GEN_2 : _T_7916_28;
  assign _GEN_195 = 5'h1d == _T_328 ? _GEN_2 : _T_7916_29;
  assign _GEN_196 = 5'h1e == _T_328 ? _GEN_2 : _T_7916_30;
  assign _GEN_197 = 5'h1f == _T_328 ? _GEN_2 : _T_7916_31;
  assign _GEN_198 = _T_7962 ? _GEN_166 : _T_7916_0;
  assign _GEN_199 = _T_7962 ? _GEN_167 : _T_7916_1;
  assign _GEN_200 = _T_7962 ? _GEN_168 : _T_7916_2;
  assign _GEN_201 = _T_7962 ? _GEN_169 : _T_7916_3;
  assign _GEN_202 = _T_7962 ? _GEN_170 : _T_7916_4;
  assign _GEN_203 = _T_7962 ? _GEN_171 : _T_7916_5;
  assign _GEN_204 = _T_7962 ? _GEN_172 : _T_7916_6;
  assign _GEN_205 = _T_7962 ? _GEN_173 : _T_7916_7;
  assign _GEN_206 = _T_7962 ? _GEN_174 : _T_7916_8;
  assign _GEN_207 = _T_7962 ? _GEN_175 : _T_7916_9;
  assign _GEN_208 = _T_7962 ? _GEN_176 : _T_7916_10;
  assign _GEN_209 = _T_7962 ? _GEN_177 : _T_7916_11;
  assign _GEN_210 = _T_7962 ? _GEN_178 : _T_7916_12;
  assign _GEN_211 = _T_7962 ? _GEN_179 : _T_7916_13;
  assign _GEN_212 = _T_7962 ? _GEN_180 : _T_7916_14;
  assign _GEN_213 = _T_7962 ? _GEN_181 : _T_7916_15;
  assign _GEN_214 = _T_7962 ? _GEN_182 : _T_7916_16;
  assign _GEN_215 = _T_7962 ? _GEN_183 : _T_7916_17;
  assign _GEN_216 = _T_7962 ? _GEN_184 : _T_7916_18;
  assign _GEN_217 = _T_7962 ? _GEN_185 : _T_7916_19;
  assign _GEN_218 = _T_7962 ? _GEN_186 : _T_7916_20;
  assign _GEN_219 = _T_7962 ? _GEN_187 : _T_7916_21;
  assign _GEN_220 = _T_7962 ? _GEN_188 : _T_7916_22;
  assign _GEN_221 = _T_7962 ? _GEN_189 : _T_7916_23;
  assign _GEN_222 = _T_7962 ? _GEN_190 : _T_7916_24;
  assign _GEN_223 = _T_7962 ? _GEN_191 : _T_7916_25;
  assign _GEN_224 = _T_7962 ? _GEN_192 : _T_7916_26;
  assign _GEN_225 = _T_7962 ? _GEN_193 : _T_7916_27;
  assign _GEN_226 = _T_7962 ? _GEN_194 : _T_7916_28;
  assign _GEN_227 = _T_7962 ? _GEN_195 : _T_7916_29;
  assign _GEN_228 = _T_7962 ? _GEN_196 : _T_7916_30;
  assign _GEN_229 = _T_7962 ? _GEN_197 : _T_7916_31;
  assign _T_7966 = _T_7901 & _T_322;
  assign _T_7968 = _T_7912 == 1'h0;
  assign _T_7969 = _T_7966 & _T_7968;
  assign _GEN_230 = _T_7969 ? 1'h1 : _T_7909;
  assign _T_7971 = _T_7909 & io_outputMemAddrReadys_0;
  assign _GEN_231 = _T_7971 ? 1'h0 : _GEN_230;
  assign _GEN_232 = _T_7971 ? 1'h1 : _T_7912;
  assign _T_7974 = {_T_7916_1,_T_7916_0};
  assign _T_7975 = {_T_7916_3,_T_7916_2};
  assign _T_7976 = {_T_7975,_T_7974};
  assign _T_7977 = {_T_7916_5,_T_7916_4};
  assign _T_7978 = {_T_7916_7,_T_7916_6};
  assign _T_7979 = {_T_7978,_T_7977};
  assign _T_7980 = {_T_7979,_T_7976};
  assign _T_7981 = {_T_7916_9,_T_7916_8};
  assign _T_7982 = {_T_7916_11,_T_7916_10};
  assign _T_7983 = {_T_7982,_T_7981};
  assign _T_7984 = {_T_7916_13,_T_7916_12};
  assign _T_7985 = {_T_7916_15,_T_7916_14};
  assign _T_7986 = {_T_7985,_T_7984};
  assign _T_7987 = {_T_7986,_T_7983};
  assign _T_7988 = {_T_7987,_T_7980};
  assign _T_7989 = {_T_7916_17,_T_7916_16};
  assign _T_7990 = {_T_7916_19,_T_7916_18};
  assign _T_7991 = {_T_7990,_T_7989};
  assign _T_7992 = {_T_7916_21,_T_7916_20};
  assign _T_7993 = {_T_7916_23,_T_7916_22};
  assign _T_7994 = {_T_7993,_T_7992};
  assign _T_7995 = {_T_7994,_T_7991};
  assign _T_7996 = {_T_7916_25,_T_7916_24};
  assign _T_7997 = {_T_7916_27,_T_7916_26};
  assign _T_7998 = {_T_7997,_T_7996};
  assign _T_7999 = {_T_7916_29,_T_7916_28};
  assign _T_8000 = {_T_7916_31,_T_7916_30};
  assign _T_8001 = {_T_8000,_T_7999};
  assign _T_8002 = {_T_8001,_T_7998};
  assign _T_8003 = {_T_8002,_T_7995};
  assign _T_8004 = {_T_8003,_T_7988};
  assign _T_8006 = _T_251 == 1'h0;
  assign _T_8008 = _T_8006 ? io_outputMemAddrReadys_0 : 1'h0;
  assign _T_8011 = io_outputMemBlockReadys_0 & _T_7953;
  assign _T_8013 = _T_8006 ? _T_8011 : 1'h0;
  assign _T_8014 = io_outputMemBlockReadys_0 & io_outputMemBlockValids_0;
  assign _T_8021 = _T_330 | _T_8011;
  assign _T_8022 = _T_7901 & _T_8021;
  assign _T_8027 = _T_251 + 1'h1;
  assign _T_8028 = _T_8027[0:0];
  assign _T_8029 = _T_8006 ? 1'h0 : _T_8028;
  assign _GEN_233 = _T_8022 ? _T_8029 : _T_251;
  assign _GEN_234 = _T_8022 ? 1'h0 : _GEN_165;
  assign _GEN_235 = _T_8022 ? 1'h0 : _GEN_164;
  assign _GEN_236 = _T_8022 ? 1'h0 : _GEN_232;
  assign _T_8037 = _T_8035 != 1'h1;
  assign _T_8039 = _T_8035 + 1'h1;
  assign _T_8040 = _T_8039[0:0];
  assign _GEN_237 = _T_8037 ? _T_8040 : _T_8035;
  assign _T_8090 = _T_8035 & _T_336;
  assign _T_8092 = _T_340 == 5'h1f;
  assign _T_8093 = _T_8090 & _T_8092;
  assign _GEN_238 = _T_8093 ? 1'h1 : _T_8087;
  assign _T_8096 = _T_8087 == 1'h0;
  assign _GEN_239 = 5'h0 == _T_340 ? _GEN_3 : _T_8050_0;
  assign _GEN_240 = 5'h1 == _T_340 ? _GEN_3 : _T_8050_1;
  assign _GEN_241 = 5'h2 == _T_340 ? _GEN_3 : _T_8050_2;
  assign _GEN_242 = 5'h3 == _T_340 ? _GEN_3 : _T_8050_3;
  assign _GEN_243 = 5'h4 == _T_340 ? _GEN_3 : _T_8050_4;
  assign _GEN_244 = 5'h5 == _T_340 ? _GEN_3 : _T_8050_5;
  assign _GEN_245 = 5'h6 == _T_340 ? _GEN_3 : _T_8050_6;
  assign _GEN_246 = 5'h7 == _T_340 ? _GEN_3 : _T_8050_7;
  assign _GEN_247 = 5'h8 == _T_340 ? _GEN_3 : _T_8050_8;
  assign _GEN_248 = 5'h9 == _T_340 ? _GEN_3 : _T_8050_9;
  assign _GEN_249 = 5'ha == _T_340 ? _GEN_3 : _T_8050_10;
  assign _GEN_250 = 5'hb == _T_340 ? _GEN_3 : _T_8050_11;
  assign _GEN_251 = 5'hc == _T_340 ? _GEN_3 : _T_8050_12;
  assign _GEN_252 = 5'hd == _T_340 ? _GEN_3 : _T_8050_13;
  assign _GEN_253 = 5'he == _T_340 ? _GEN_3 : _T_8050_14;
  assign _GEN_254 = 5'hf == _T_340 ? _GEN_3 : _T_8050_15;
  assign _GEN_255 = 5'h10 == _T_340 ? _GEN_3 : _T_8050_16;
  assign _GEN_256 = 5'h11 == _T_340 ? _GEN_3 : _T_8050_17;
  assign _GEN_257 = 5'h12 == _T_340 ? _GEN_3 : _T_8050_18;
  assign _GEN_258 = 5'h13 == _T_340 ? _GEN_3 : _T_8050_19;
  assign _GEN_259 = 5'h14 == _T_340 ? _GEN_3 : _T_8050_20;
  assign _GEN_260 = 5'h15 == _T_340 ? _GEN_3 : _T_8050_21;
  assign _GEN_261 = 5'h16 == _T_340 ? _GEN_3 : _T_8050_22;
  assign _GEN_262 = 5'h17 == _T_340 ? _GEN_3 : _T_8050_23;
  assign _GEN_263 = 5'h18 == _T_340 ? _GEN_3 : _T_8050_24;
  assign _GEN_264 = 5'h19 == _T_340 ? _GEN_3 : _T_8050_25;
  assign _GEN_265 = 5'h1a == _T_340 ? _GEN_3 : _T_8050_26;
  assign _GEN_266 = 5'h1b == _T_340 ? _GEN_3 : _T_8050_27;
  assign _GEN_267 = 5'h1c == _T_340 ? _GEN_3 : _T_8050_28;
  assign _GEN_268 = 5'h1d == _T_340 ? _GEN_3 : _T_8050_29;
  assign _GEN_269 = 5'h1e == _T_340 ? _GEN_3 : _T_8050_30;
  assign _GEN_270 = 5'h1f == _T_340 ? _GEN_3 : _T_8050_31;
  assign _GEN_271 = _T_8096 ? _GEN_239 : _T_8050_0;
  assign _GEN_272 = _T_8096 ? _GEN_240 : _T_8050_1;
  assign _GEN_273 = _T_8096 ? _GEN_241 : _T_8050_2;
  assign _GEN_274 = _T_8096 ? _GEN_242 : _T_8050_3;
  assign _GEN_275 = _T_8096 ? _GEN_243 : _T_8050_4;
  assign _GEN_276 = _T_8096 ? _GEN_244 : _T_8050_5;
  assign _GEN_277 = _T_8096 ? _GEN_245 : _T_8050_6;
  assign _GEN_278 = _T_8096 ? _GEN_246 : _T_8050_7;
  assign _GEN_279 = _T_8096 ? _GEN_247 : _T_8050_8;
  assign _GEN_280 = _T_8096 ? _GEN_248 : _T_8050_9;
  assign _GEN_281 = _T_8096 ? _GEN_249 : _T_8050_10;
  assign _GEN_282 = _T_8096 ? _GEN_250 : _T_8050_11;
  assign _GEN_283 = _T_8096 ? _GEN_251 : _T_8050_12;
  assign _GEN_284 = _T_8096 ? _GEN_252 : _T_8050_13;
  assign _GEN_285 = _T_8096 ? _GEN_253 : _T_8050_14;
  assign _GEN_286 = _T_8096 ? _GEN_254 : _T_8050_15;
  assign _GEN_287 = _T_8096 ? _GEN_255 : _T_8050_16;
  assign _GEN_288 = _T_8096 ? _GEN_256 : _T_8050_17;
  assign _GEN_289 = _T_8096 ? _GEN_257 : _T_8050_18;
  assign _GEN_290 = _T_8096 ? _GEN_258 : _T_8050_19;
  assign _GEN_291 = _T_8096 ? _GEN_259 : _T_8050_20;
  assign _GEN_292 = _T_8096 ? _GEN_260 : _T_8050_21;
  assign _GEN_293 = _T_8096 ? _GEN_261 : _T_8050_22;
  assign _GEN_294 = _T_8096 ? _GEN_262 : _T_8050_23;
  assign _GEN_295 = _T_8096 ? _GEN_263 : _T_8050_24;
  assign _GEN_296 = _T_8096 ? _GEN_264 : _T_8050_25;
  assign _GEN_297 = _T_8096 ? _GEN_265 : _T_8050_26;
  assign _GEN_298 = _T_8096 ? _GEN_266 : _T_8050_27;
  assign _GEN_299 = _T_8096 ? _GEN_267 : _T_8050_28;
  assign _GEN_300 = _T_8096 ? _GEN_268 : _T_8050_29;
  assign _GEN_301 = _T_8096 ? _GEN_269 : _T_8050_30;
  assign _GEN_302 = _T_8096 ? _GEN_270 : _T_8050_31;
  assign _T_8100 = _T_8035 & _T_334;
  assign _T_8102 = _T_8046 == 1'h0;
  assign _T_8103 = _T_8100 & _T_8102;
  assign _GEN_303 = _T_8103 ? 1'h1 : _T_8043;
  assign _T_8105 = _T_8043 & io_outputMemAddrReadys_1;
  assign _GEN_304 = _T_8105 ? 1'h0 : _GEN_303;
  assign _GEN_305 = _T_8105 ? 1'h1 : _T_8046;
  assign _T_8108 = {_T_8050_1,_T_8050_0};
  assign _T_8109 = {_T_8050_3,_T_8050_2};
  assign _T_8110 = {_T_8109,_T_8108};
  assign _T_8111 = {_T_8050_5,_T_8050_4};
  assign _T_8112 = {_T_8050_7,_T_8050_6};
  assign _T_8113 = {_T_8112,_T_8111};
  assign _T_8114 = {_T_8113,_T_8110};
  assign _T_8115 = {_T_8050_9,_T_8050_8};
  assign _T_8116 = {_T_8050_11,_T_8050_10};
  assign _T_8117 = {_T_8116,_T_8115};
  assign _T_8118 = {_T_8050_13,_T_8050_12};
  assign _T_8119 = {_T_8050_15,_T_8050_14};
  assign _T_8120 = {_T_8119,_T_8118};
  assign _T_8121 = {_T_8120,_T_8117};
  assign _T_8122 = {_T_8121,_T_8114};
  assign _T_8123 = {_T_8050_17,_T_8050_16};
  assign _T_8124 = {_T_8050_19,_T_8050_18};
  assign _T_8125 = {_T_8124,_T_8123};
  assign _T_8126 = {_T_8050_21,_T_8050_20};
  assign _T_8127 = {_T_8050_23,_T_8050_22};
  assign _T_8128 = {_T_8127,_T_8126};
  assign _T_8129 = {_T_8128,_T_8125};
  assign _T_8130 = {_T_8050_25,_T_8050_24};
  assign _T_8131 = {_T_8050_27,_T_8050_26};
  assign _T_8132 = {_T_8131,_T_8130};
  assign _T_8133 = {_T_8050_29,_T_8050_28};
  assign _T_8134 = {_T_8050_31,_T_8050_30};
  assign _T_8135 = {_T_8134,_T_8133};
  assign _T_8136 = {_T_8135,_T_8132};
  assign _T_8137 = {_T_8136,_T_8129};
  assign _T_8138 = {_T_8137,_T_8122};
  assign _T_8142 = _T_254 ? io_outputMemAddrReadys_1 : 1'h0;
  assign _T_8145 = io_outputMemBlockReadys_1 & _T_8087;
  assign _T_8147 = _T_254 ? _T_8145 : 1'h0;
  assign _T_8148 = io_outputMemBlockReadys_1 & io_outputMemBlockValids_1;
  assign _T_8155 = _T_342 | _T_8145;
  assign _T_8156 = _T_8035 & _T_8155;
  assign _T_8161 = _T_254 + 1'h1;
  assign _T_8162 = _T_8161[0:0];
  assign _T_8163 = _T_254 ? 1'h1 : _T_8162;
  assign _GEN_306 = _T_8156 ? _T_8163 : _T_254;
  assign _GEN_307 = _T_8156 ? 1'h0 : _GEN_238;
  assign _GEN_308 = _T_8156 ? 1'h0 : _GEN_237;
  assign _GEN_309 = _T_8156 ? 1'h0 : _GEN_305;
  assign cumFinished = cores_0_outputFinished & cores_1_outputFinished;
  assign io_inputMemAddrs_0 = _T_265_0;
  assign io_inputMemAddrs_1 = _T_297_0;
  assign io_inputMemAddrValids_0 = _T_382;
  assign io_inputMemAddrValids_1 = _T_4160;
  assign io_inputMemBlockReadys_0 = _T_4106;
  assign io_inputMemBlockReadys_1 = _T_7884;
  assign io_outputMemAddrs_0 = _T_320;
  assign io_outputMemAddrs_1 = _T_332;
  assign io_outputMemAddrValids_0 = _T_7909;
  assign io_outputMemAddrValids_1 = _T_8043;
  assign io_outputMemBlocks_0 = _T_8004;
  assign io_outputMemBlocks_1 = _T_8138;
  assign io_outputMemBlockValids_0 = _T_7953;
  assign io_outputMemBlockValids_1 = _T_8087;
  assign io_finished = cumFinished;
  assign StreamingCore_io_inputMemAddrConsumed = cores_0_inputMemAddrConsumed;
  assign StreamingCore_io_inputMemBlock = cores_0_inputMemBlock;
  assign StreamingCore_io_inputMemIdx = cores_0_inputMemIdx;
  assign StreamingCore_io_inputMemBlockValid = cores_0_inputMemBlockValid;
  assign StreamingCore_io_outputMemAddrReady = cores_0_outputMemAddrReady;
  assign StreamingCore_io_outputMemBlockReady = cores_0_outputMemBlockReady;
  assign StreamingCore_clock = clock;
  assign StreamingCore_reset = reset;
  assign StreamingCore_1_io_inputMemAddrConsumed = cores_1_inputMemAddrConsumed;
  assign StreamingCore_1_io_inputMemBlock = cores_1_inputMemBlock;
  assign StreamingCore_1_io_inputMemIdx = cores_1_inputMemIdx;
  assign StreamingCore_1_io_inputMemBlockValid = cores_1_inputMemBlockValid;
  assign StreamingCore_1_io_outputMemAddrReady = cores_1_outputMemAddrReady;
  assign StreamingCore_1_io_outputMemBlockReady = cores_1_outputMemBlockReady;
  assign StreamingCore_1_clock = clock;
  assign StreamingCore_1_reset = reset;
  assign cores_0_inputMemAddr = StreamingCore_io_inputMemAddr;
  assign cores_0_inputMemAddrConsumed = _T_4114;
  assign cores_0_inputMemBlock = _GEN_0;
  assign cores_0_inputMemIdx = _T_683_0;
  assign cores_0_inputMemBlockValid = _T_4120;
  assign cores_0_inputMemBlockReady = StreamingCore_io_inputMemBlockReady;
  assign cores_0_outputMemAddr = StreamingCore_io_outputMemAddr;
  assign cores_0_outputMemAddrValid = StreamingCore_io_outputMemAddrValid;
  assign cores_0_outputMemAddrReady = _T_8008;
  assign cores_0_outputMemBlock = StreamingCore_io_outputMemBlock;
  assign cores_0_outputMemIdx = StreamingCore_io_outputMemIdx;
  assign cores_0_outputMemBlockValid = StreamingCore_io_outputMemBlockValid;
  assign cores_0_outputMemBlockReady = _T_8013;
  assign cores_0_inputAddrsIgnore = StreamingCore_io_inputAddrsIgnore;
  assign cores_0_inputBlocksFinished = StreamingCore_io_inputBlocksFinished;
  assign cores_0_outputFinished = StreamingCore_io_outputFinished;
  assign cores_1_inputMemAddr = StreamingCore_1_io_inputMemAddr;
  assign cores_1_inputMemAddrConsumed = _T_7892;
  assign cores_1_inputMemBlock = _GEN_1;
  assign cores_1_inputMemIdx = _T_4461_0;
  assign cores_1_inputMemBlockValid = _T_7898;
  assign cores_1_inputMemBlockReady = StreamingCore_1_io_inputMemBlockReady;
  assign cores_1_outputMemAddr = StreamingCore_1_io_outputMemAddr;
  assign cores_1_outputMemAddrValid = StreamingCore_1_io_outputMemAddrValid;
  assign cores_1_outputMemAddrReady = _T_8142;
  assign cores_1_outputMemBlock = StreamingCore_1_io_outputMemBlock;
  assign cores_1_outputMemIdx = StreamingCore_1_io_outputMemIdx;
  assign cores_1_outputMemBlockValid = StreamingCore_1_io_outputMemBlockValid;
  assign cores_1_outputMemBlockReady = _T_8147;
  assign cores_1_inputAddrsIgnore = StreamingCore_1_io_inputAddrsIgnore;
  assign cores_1_inputBlocksFinished = StreamingCore_1_io_inputBlocksFinished;
  assign cores_1_outputFinished = StreamingCore_1_io_outputFinished;
  assign _T_265_0 = _T_256;
  assign _T_271_0 = _T_258;
  assign _T_277_0 = _T_260;
  assign _T_283_0 = _T_262;
  assign _T_297_0 = _T_288;
  assign _T_303_0 = _T_290;
  assign _T_309_0 = _T_292;
  assign _T_315_0 = _T_294;
  assign _GEN_0 = _GEN_83;
  assign _GEN_1 = _GEN_163;
  assign _GEN_2 = _T_326;
  assign _GEN_3 = _T_338;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_239 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_242 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_245 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_248 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_251 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_254 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{$random}};
  _T_256 = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_258 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_260 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_262 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{$random}};
  _T_288 = _RAND_10[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_290 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_292 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_294 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{$random}};
  _T_320 = _RAND_14[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_322 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_324 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_326 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_328 = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_330 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{$random}};
  _T_332 = _RAND_20[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_334 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_336 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_338 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_340 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_342 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_345 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_353 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_385 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_464_0_0 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_464_0_1 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_464_0_2 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_464_0_3 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_464_0_4 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_464_0_5 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_464_0_6 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_464_0_7 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_464_0_8 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_464_0_9 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_464_0_10 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_464_0_11 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_464_0_12 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_464_0_13 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_464_0_14 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_464_0_15 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_464_0_16 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_464_0_17 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_464_0_18 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_464_0_19 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_464_0_20 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_464_0_21 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_464_0_22 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_464_0_23 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_464_0_24 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_464_0_25 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_464_0_26 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_464_0_27 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_464_0_28 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_464_0_29 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_464_0_30 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_464_0_31 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_683_0 = _RAND_61[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_704_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_714 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_4123 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_4131 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_4163 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_4242_0_0 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_4242_0_1 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_4242_0_2 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_4242_0_3 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_4242_0_4 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_4242_0_5 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_4242_0_6 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_4242_0_7 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_4242_0_8 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_4242_0_9 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_4242_0_10 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_4242_0_11 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_4242_0_12 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_4242_0_13 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_4242_0_14 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_4242_0_15 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_4242_0_16 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_4242_0_17 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_4242_0_18 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_4242_0_19 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_4242_0_20 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_4242_0_21 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_4242_0_22 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_4242_0_23 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_4242_0_24 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_4242_0_25 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_4242_0_26 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_4242_0_27 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_4242_0_28 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_4242_0_29 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_4242_0_30 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_4242_0_31 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_4461_0 = _RAND_99[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_4482_0 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_4492 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_7901 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_7909 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_7912 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_7916_0 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_7916_1 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_7916_2 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_7916_3 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_7916_4 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_7916_5 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_7916_6 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_7916_7 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_7916_8 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_7916_9 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_7916_10 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_7916_11 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_7916_12 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_7916_13 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_7916_14 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_7916_15 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_7916_16 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_7916_17 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_7916_18 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_7916_19 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_7916_20 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_7916_21 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_7916_22 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_7916_23 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_7916_24 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_7916_25 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_7916_26 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_7916_27 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_7916_28 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_7916_29 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  _T_7916_30 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_7916_31 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  _T_7953 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  _T_8035 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  _T_8043 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  _T_8046 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  _T_8050_0 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  _T_8050_1 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  _T_8050_2 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  _T_8050_3 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  _T_8050_4 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  _T_8050_5 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  _T_8050_6 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  _T_8050_7 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  _T_8050_8 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  _T_8050_9 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  _T_8050_10 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  _T_8050_11 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  _T_8050_12 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  _T_8050_13 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _T_8050_14 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  _T_8050_15 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _T_8050_16 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  _T_8050_17 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  _T_8050_18 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _T_8050_19 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  _T_8050_20 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  _T_8050_21 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  _T_8050_22 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  _T_8050_23 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  _T_8050_24 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  _T_8050_25 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  _T_8050_26 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  _T_8050_27 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  _T_8050_28 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  _T_8050_29 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  _T_8050_30 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  _T_8050_31 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  _T_8087 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      if (_T_359) begin
        if (_T_361) begin
          if (_T_363) begin
            _T_239 <= 1'h0;
          end else begin
            _T_239 <= _T_367;
          end
        end
      end
    end
    if (reset) begin
      _T_242 <= 1'h0;
    end else begin
      if (_T_4070) begin
        if (_T_4072) begin
          _T_242 <= 1'h0;
        end else begin
          _T_242 <= _T_4076;
        end
      end
    end
    if (reset) begin
      _T_245 <= 1'h1;
    end else begin
      if (_T_4137) begin
        if (_T_4139) begin
          if (_T_245) begin
            _T_245 <= 1'h1;
          end else begin
            _T_245 <= _T_4145;
          end
        end
      end
    end
    if (reset) begin
      _T_248 <= 1'h1;
    end else begin
      if (_T_7848) begin
        if (_T_248) begin
          _T_248 <= 1'h1;
        end else begin
          _T_248 <= _T_7854;
        end
      end
    end
    if (reset) begin
      _T_251 <= 1'h0;
    end else begin
      if (_T_8022) begin
        if (_T_8006) begin
          _T_251 <= 1'h0;
        end else begin
          _T_251 <= _T_8028;
        end
      end
    end
    if (reset) begin
      _T_254 <= 1'h1;
    end else begin
      if (_T_8156) begin
        if (_T_254) begin
          _T_254 <= 1'h1;
        end else begin
          _T_254 <= _T_8162;
        end
      end
    end
    _T_256 <= {{32'd0}, cores_0_inputMemAddr};
    _T_258 <= cores_0_inputMemBlockReady;
    _T_260 <= cores_0_inputAddrsIgnore;
    _T_262 <= cores_0_inputBlocksFinished;
    _T_288 <= {{32'd0}, cores_1_inputMemAddr};
    _T_290 <= cores_1_inputMemBlockReady;
    _T_292 <= cores_1_inputAddrsIgnore;
    _T_294 <= cores_1_inputBlocksFinished;
    _T_320 <= {{32'd0}, cores_0_outputMemAddr};
    _T_322 <= cores_0_outputMemAddrValid;
    _T_324 <= cores_0_outputMemBlockValid;
    _T_326 <= cores_0_outputMemBlock;
    _T_328 <= cores_0_outputMemIdx;
    _T_330 <= cores_0_outputFinished;
    _T_332 <= {{32'd0}, cores_1_outputMemAddr};
    _T_334 <= cores_1_outputMemAddrValid;
    _T_336 <= cores_1_outputMemBlockValid;
    _T_338 <= cores_1_outputMemBlock;
    _T_340 <= cores_1_outputMemIdx;
    _T_342 <= cores_1_outputFinished;
    if (reset) begin
      _T_345 <= 1'h0;
    end else begin
      if (_T_359) begin
        if (_T_361) begin
          _T_345 <= 1'h0;
        end else begin
          if (_T_347) begin
            _T_345 <= _T_350;
          end
        end
      end else begin
        if (_T_347) begin
          _T_345 <= _T_350;
        end
      end
    end
    if (reset) begin
      _T_353 <= 1'h0;
    end else begin
      if (_T_359) begin
        if (_T_361) begin
          _T_353 <= 1'h0;
        end else begin
          _T_353 <= _T_373;
        end
      end
    end
    if (reset) begin
      _T_385 <= 1'h0;
    end else begin
      if (_T_4070) begin
        _T_385 <= 1'h0;
      end else begin
        if (_T_387) begin
          _T_385 <= _T_390;
        end
      end
    end
    if (_T_726) begin
      _T_464_0_0 <= _T_830;
    end
    if (_T_726) begin
      _T_464_0_1 <= _T_934;
    end
    if (_T_726) begin
      _T_464_0_2 <= _T_1038;
    end
    if (_T_726) begin
      _T_464_0_3 <= _T_1142;
    end
    if (_T_726) begin
      _T_464_0_4 <= _T_1246;
    end
    if (_T_726) begin
      _T_464_0_5 <= _T_1350;
    end
    if (_T_726) begin
      _T_464_0_6 <= _T_1454;
    end
    if (_T_726) begin
      _T_464_0_7 <= _T_1558;
    end
    if (_T_726) begin
      _T_464_0_8 <= _T_1662;
    end
    if (_T_726) begin
      _T_464_0_9 <= _T_1766;
    end
    if (_T_726) begin
      _T_464_0_10 <= _T_1870;
    end
    if (_T_726) begin
      _T_464_0_11 <= _T_1974;
    end
    if (_T_726) begin
      _T_464_0_12 <= _T_2078;
    end
    if (_T_726) begin
      _T_464_0_13 <= _T_2182;
    end
    if (_T_726) begin
      _T_464_0_14 <= _T_2286;
    end
    if (_T_726) begin
      _T_464_0_15 <= _T_2390;
    end
    if (_T_726) begin
      _T_464_0_16 <= _T_2494;
    end
    if (_T_726) begin
      _T_464_0_17 <= _T_2598;
    end
    if (_T_726) begin
      _T_464_0_18 <= _T_2702;
    end
    if (_T_726) begin
      _T_464_0_19 <= _T_2806;
    end
    if (_T_726) begin
      _T_464_0_20 <= _T_2910;
    end
    if (_T_726) begin
      _T_464_0_21 <= _T_3014;
    end
    if (_T_726) begin
      _T_464_0_22 <= _T_3118;
    end
    if (_T_726) begin
      _T_464_0_23 <= _T_3222;
    end
    if (_T_726) begin
      _T_464_0_24 <= _T_3326;
    end
    if (_T_726) begin
      _T_464_0_25 <= _T_3430;
    end
    if (_T_726) begin
      _T_464_0_26 <= _T_3534;
    end
    if (_T_726) begin
      _T_464_0_27 <= _T_3638;
    end
    if (_T_726) begin
      _T_464_0_28 <= _T_3742;
    end
    if (_T_726) begin
      _T_464_0_29 <= _T_3846;
    end
    if (_T_726) begin
      _T_464_0_30 <= _T_3950;
    end
    if (_T_726) begin
      _T_464_0_31 <= _T_4054;
    end
    if (reset) begin
      _T_683_0 <= 5'h0;
    end else begin
      if (_T_704_0) begin
        if (_T_4086) begin
          _T_683_0 <= 5'h0;
        end else begin
          _T_683_0 <= _T_4091;
        end
      end
    end
    if (reset) begin
      _T_704_0 <= 1'h0;
    end else begin
      if (_T_704_0) begin
        if (_T_4086) begin
          _T_704_0 <= 1'h0;
        end else begin
          if (_T_726) begin
            _T_704_0 <= _T_4062;
          end
        end
      end else begin
        if (_T_726) begin
          _T_704_0 <= _T_4062;
        end
      end
    end
    if (reset) begin
      _T_714 <= 1'h0;
    end else begin
      if (_T_4070) begin
        _T_714 <= 1'h0;
      end else begin
        if (_T_726) begin
          _T_714 <= _T_4065;
        end
      end
    end
    if (reset) begin
      _T_4123 <= 1'h0;
    end else begin
      if (_T_4137) begin
        if (_T_4139) begin
          _T_4123 <= 1'h0;
        end else begin
          if (_T_4125) begin
            _T_4123 <= _T_4128;
          end
        end
      end else begin
        if (_T_4125) begin
          _T_4123 <= _T_4128;
        end
      end
    end
    if (reset) begin
      _T_4131 <= 1'h0;
    end else begin
      if (_T_4137) begin
        if (_T_4139) begin
          _T_4131 <= 1'h0;
        end else begin
          _T_4131 <= _T_4151;
        end
      end
    end
    if (reset) begin
      _T_4163 <= 1'h0;
    end else begin
      if (_T_7848) begin
        _T_4163 <= 1'h0;
      end else begin
        if (_T_4165) begin
          _T_4163 <= _T_4168;
        end
      end
    end
    if (_T_4504) begin
      _T_4242_0_0 <= _T_4608;
    end
    if (_T_4504) begin
      _T_4242_0_1 <= _T_4712;
    end
    if (_T_4504) begin
      _T_4242_0_2 <= _T_4816;
    end
    if (_T_4504) begin
      _T_4242_0_3 <= _T_4920;
    end
    if (_T_4504) begin
      _T_4242_0_4 <= _T_5024;
    end
    if (_T_4504) begin
      _T_4242_0_5 <= _T_5128;
    end
    if (_T_4504) begin
      _T_4242_0_6 <= _T_5232;
    end
    if (_T_4504) begin
      _T_4242_0_7 <= _T_5336;
    end
    if (_T_4504) begin
      _T_4242_0_8 <= _T_5440;
    end
    if (_T_4504) begin
      _T_4242_0_9 <= _T_5544;
    end
    if (_T_4504) begin
      _T_4242_0_10 <= _T_5648;
    end
    if (_T_4504) begin
      _T_4242_0_11 <= _T_5752;
    end
    if (_T_4504) begin
      _T_4242_0_12 <= _T_5856;
    end
    if (_T_4504) begin
      _T_4242_0_13 <= _T_5960;
    end
    if (_T_4504) begin
      _T_4242_0_14 <= _T_6064;
    end
    if (_T_4504) begin
      _T_4242_0_15 <= _T_6168;
    end
    if (_T_4504) begin
      _T_4242_0_16 <= _T_6272;
    end
    if (_T_4504) begin
      _T_4242_0_17 <= _T_6376;
    end
    if (_T_4504) begin
      _T_4242_0_18 <= _T_6480;
    end
    if (_T_4504) begin
      _T_4242_0_19 <= _T_6584;
    end
    if (_T_4504) begin
      _T_4242_0_20 <= _T_6688;
    end
    if (_T_4504) begin
      _T_4242_0_21 <= _T_6792;
    end
    if (_T_4504) begin
      _T_4242_0_22 <= _T_6896;
    end
    if (_T_4504) begin
      _T_4242_0_23 <= _T_7000;
    end
    if (_T_4504) begin
      _T_4242_0_24 <= _T_7104;
    end
    if (_T_4504) begin
      _T_4242_0_25 <= _T_7208;
    end
    if (_T_4504) begin
      _T_4242_0_26 <= _T_7312;
    end
    if (_T_4504) begin
      _T_4242_0_27 <= _T_7416;
    end
    if (_T_4504) begin
      _T_4242_0_28 <= _T_7520;
    end
    if (_T_4504) begin
      _T_4242_0_29 <= _T_7624;
    end
    if (_T_4504) begin
      _T_4242_0_30 <= _T_7728;
    end
    if (_T_4504) begin
      _T_4242_0_31 <= _T_7832;
    end
    if (reset) begin
      _T_4461_0 <= 5'h0;
    end else begin
      if (_T_4482_0) begin
        if (_T_7864) begin
          _T_4461_0 <= 5'h0;
        end else begin
          _T_4461_0 <= _T_7869;
        end
      end
    end
    if (reset) begin
      _T_4482_0 <= 1'h0;
    end else begin
      if (_T_4482_0) begin
        if (_T_7864) begin
          _T_4482_0 <= 1'h0;
        end else begin
          if (_T_4504) begin
            _T_4482_0 <= _T_7840;
          end
        end
      end else begin
        if (_T_4504) begin
          _T_4482_0 <= _T_7840;
        end
      end
    end
    if (reset) begin
      _T_4492 <= 1'h0;
    end else begin
      if (_T_7848) begin
        _T_4492 <= 1'h0;
      end else begin
        if (_T_4504) begin
          _T_4492 <= _T_7843;
        end
      end
    end
    if (reset) begin
      _T_7901 <= 1'h0;
    end else begin
      if (_T_8022) begin
        _T_7901 <= 1'h0;
      end else begin
        if (_T_7903) begin
          _T_7901 <= _T_7906;
        end
      end
    end
    if (reset) begin
      _T_7909 <= 1'h0;
    end else begin
      if (_T_7971) begin
        _T_7909 <= 1'h0;
      end else begin
        if (_T_7969) begin
          _T_7909 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_7912 <= 1'h0;
    end else begin
      if (_T_8022) begin
        _T_7912 <= 1'h0;
      end else begin
        if (_T_7971) begin
          _T_7912 <= 1'h1;
        end
      end
    end
    if (_T_7962) begin
      if (5'h0 == _T_328) begin
        _T_7916_0 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h1 == _T_328) begin
        _T_7916_1 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h2 == _T_328) begin
        _T_7916_2 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h3 == _T_328) begin
        _T_7916_3 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h4 == _T_328) begin
        _T_7916_4 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h5 == _T_328) begin
        _T_7916_5 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h6 == _T_328) begin
        _T_7916_6 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h7 == _T_328) begin
        _T_7916_7 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h8 == _T_328) begin
        _T_7916_8 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h9 == _T_328) begin
        _T_7916_9 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'ha == _T_328) begin
        _T_7916_10 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'hb == _T_328) begin
        _T_7916_11 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'hc == _T_328) begin
        _T_7916_12 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'hd == _T_328) begin
        _T_7916_13 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'he == _T_328) begin
        _T_7916_14 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'hf == _T_328) begin
        _T_7916_15 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h10 == _T_328) begin
        _T_7916_16 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h11 == _T_328) begin
        _T_7916_17 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h12 == _T_328) begin
        _T_7916_18 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h13 == _T_328) begin
        _T_7916_19 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h14 == _T_328) begin
        _T_7916_20 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h15 == _T_328) begin
        _T_7916_21 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h16 == _T_328) begin
        _T_7916_22 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h17 == _T_328) begin
        _T_7916_23 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h18 == _T_328) begin
        _T_7916_24 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h19 == _T_328) begin
        _T_7916_25 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h1a == _T_328) begin
        _T_7916_26 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h1b == _T_328) begin
        _T_7916_27 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h1c == _T_328) begin
        _T_7916_28 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h1d == _T_328) begin
        _T_7916_29 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h1e == _T_328) begin
        _T_7916_30 <= _GEN_2;
      end
    end
    if (_T_7962) begin
      if (5'h1f == _T_328) begin
        _T_7916_31 <= _GEN_2;
      end
    end
    if (reset) begin
      _T_7953 <= 1'h0;
    end else begin
      if (_T_8022) begin
        _T_7953 <= 1'h0;
      end else begin
        if (_T_7959) begin
          _T_7953 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_8035 <= 1'h0;
    end else begin
      if (_T_8156) begin
        _T_8035 <= 1'h0;
      end else begin
        if (_T_8037) begin
          _T_8035 <= _T_8040;
        end
      end
    end
    if (reset) begin
      _T_8043 <= 1'h0;
    end else begin
      if (_T_8105) begin
        _T_8043 <= 1'h0;
      end else begin
        if (_T_8103) begin
          _T_8043 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_8046 <= 1'h0;
    end else begin
      if (_T_8156) begin
        _T_8046 <= 1'h0;
      end else begin
        if (_T_8105) begin
          _T_8046 <= 1'h1;
        end
      end
    end
    if (_T_8096) begin
      if (5'h0 == _T_340) begin
        _T_8050_0 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h1 == _T_340) begin
        _T_8050_1 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h2 == _T_340) begin
        _T_8050_2 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h3 == _T_340) begin
        _T_8050_3 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h4 == _T_340) begin
        _T_8050_4 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h5 == _T_340) begin
        _T_8050_5 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h6 == _T_340) begin
        _T_8050_6 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h7 == _T_340) begin
        _T_8050_7 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h8 == _T_340) begin
        _T_8050_8 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h9 == _T_340) begin
        _T_8050_9 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'ha == _T_340) begin
        _T_8050_10 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'hb == _T_340) begin
        _T_8050_11 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'hc == _T_340) begin
        _T_8050_12 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'hd == _T_340) begin
        _T_8050_13 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'he == _T_340) begin
        _T_8050_14 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'hf == _T_340) begin
        _T_8050_15 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h10 == _T_340) begin
        _T_8050_16 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h11 == _T_340) begin
        _T_8050_17 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h12 == _T_340) begin
        _T_8050_18 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h13 == _T_340) begin
        _T_8050_19 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h14 == _T_340) begin
        _T_8050_20 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h15 == _T_340) begin
        _T_8050_21 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h16 == _T_340) begin
        _T_8050_22 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h17 == _T_340) begin
        _T_8050_23 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h18 == _T_340) begin
        _T_8050_24 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h19 == _T_340) begin
        _T_8050_25 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h1a == _T_340) begin
        _T_8050_26 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h1b == _T_340) begin
        _T_8050_27 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h1c == _T_340) begin
        _T_8050_28 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h1d == _T_340) begin
        _T_8050_29 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h1e == _T_340) begin
        _T_8050_30 <= _GEN_3;
      end
    end
    if (_T_8096) begin
      if (5'h1f == _T_340) begin
        _T_8050_31 <= _GEN_3;
      end
    end
    if (reset) begin
      _T_8087 <= 1'h0;
    end else begin
      if (_T_8156) begin
        _T_8087 <= 1'h0;
      end else begin
        if (_T_8093) begin
          _T_8087 <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_722 & _T_4084) begin
          $fwrite(32'h80000002,"inputBuffer: 0x%h for core %d, channel 0\n",io_inputMemBlocks_0,_T_4081);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4500 & _T_4084) begin
          $fwrite(32'h80000002,"inputBuffer: 0x%h for core %d, channel 1\n",io_inputMemBlocks_1,_T_7859);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8014 & _T_4084) begin
          $fwrite(32'h80000002,"outputBuffer: 0x%h for core %d, channel 0\n",io_outputMemBlocks_0,_T_251);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8148 & _T_4084) begin
          $fwrite(32'h80000002,"outputBuffer: 0x%h for core %d, channel 1\n",io_outputMemBlocks_1,_T_254);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
