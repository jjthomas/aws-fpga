`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module DualPortBRAM(
  input         clock,
  input  [4:0]  io_a_addr,
  input  [15:0] io_a_din,
  input         io_a_wr,
  input  [4:0]  io_b_addr,
  output [15:0] io_b_dout
);
  reg [15:0] mem [0:31];
  reg [31:0] _RAND_0;
  wire [15:0] mem__T_12_data;
  wire [4:0] mem__T_12_addr;
  wire [15:0] mem__T_14_data;
  wire [4:0] mem__T_14_addr;
  wire [15:0] mem__T_13_data;
  wire [4:0] mem__T_13_addr;
  wire  mem__T_13_mask;
  wire  mem__T_13_en;
  wire [15:0] mem__T_15_data;
  wire [4:0] mem__T_15_addr;
  wire  mem__T_15_mask;
  wire  mem__T_15_en;
  wire  _GEN_8;
  reg [4:0] mem__T_12_addr_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] mem__T_14_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign mem__T_12_addr = mem__T_12_addr_pipe_0;
  assign mem__T_12_data = mem[mem__T_12_addr];
  assign mem__T_14_addr = mem__T_14_addr_pipe_0;
  assign mem__T_14_data = mem[mem__T_14_addr];
  assign mem__T_13_data = io_a_din;
  assign mem__T_13_addr = io_a_addr;
  assign mem__T_13_mask = io_a_wr;
  assign mem__T_13_en = io_a_wr;
  assign mem__T_15_data = 16'h0;
  assign mem__T_15_addr = io_b_addr;
  assign mem__T_15_mask = 1'h0;
  assign mem__T_15_en = 1'h0;
  assign _GEN_8 = 1'h1;
  assign io_b_dout = mem__T_14_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem__T_12_addr_pipe_0 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem__T_14_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_13_en & mem__T_13_mask) begin
      mem[mem__T_13_addr] <= mem__T_13_data;
    end
    if(mem__T_15_en & mem__T_15_mask) begin
      mem[mem__T_15_addr] <= mem__T_15_data;
    end
    if (_GEN_8) begin
      mem__T_12_addr_pipe_0 <= io_a_addr;
    end
    if (_GEN_8) begin
      mem__T_14_addr_pipe_0 <= io_b_addr;
    end
  end
endmodule
module PassThrough(
  input         clock,
  input         reset,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  input  [9:0]  io_inputBits,
  output        io_inputMemConsumed,
  input         io_inputFinished,
  output [15:0] io_outputMemBlock,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output [9:0]  io_outputBits,
  output        io_outputFinished,
  input         io_outputMemFlushed
);
  reg  inputMemBlock_0;
  reg [31:0] _RAND_0;
  reg  inputMemBlock_1;
  reg [31:0] _RAND_1;
  reg  inputMemBlock_2;
  reg [31:0] _RAND_2;
  reg  inputMemBlock_3;
  reg [31:0] _RAND_3;
  reg  inputMemBlock_4;
  reg [31:0] _RAND_4;
  reg  inputMemBlock_5;
  reg [31:0] _RAND_5;
  reg  inputMemBlock_6;
  reg [31:0] _RAND_6;
  reg  inputMemBlock_7;
  reg [31:0] _RAND_7;
  reg  inputMemBlock_8;
  reg [31:0] _RAND_8;
  reg  inputMemBlock_9;
  reg [31:0] _RAND_9;
  reg  inputMemBlock_10;
  reg [31:0] _RAND_10;
  reg  inputMemBlock_11;
  reg [31:0] _RAND_11;
  reg  inputMemBlock_12;
  reg [31:0] _RAND_12;
  reg  inputMemBlock_13;
  reg [31:0] _RAND_13;
  reg  inputMemBlock_14;
  reg [31:0] _RAND_14;
  reg  inputMemBlock_15;
  reg [31:0] _RAND_15;
  reg [4:0] inputPieceBitsRemaining;
  reg [31:0] _RAND_16;
  reg [9:0] inputBitsRemaining;
  reg [31:0] _RAND_17;
  reg  inputBlockLoaded;
  reg [31:0] _RAND_18;
  reg  outputMemBlock_0;
  reg [31:0] _RAND_19;
  reg  outputMemBlock_1;
  reg [31:0] _RAND_20;
  reg  outputMemBlock_2;
  reg [31:0] _RAND_21;
  reg  outputMemBlock_3;
  reg [31:0] _RAND_22;
  reg  outputMemBlock_4;
  reg [31:0] _RAND_23;
  reg  outputMemBlock_5;
  reg [31:0] _RAND_24;
  reg  outputMemBlock_6;
  reg [31:0] _RAND_25;
  reg  outputMemBlock_7;
  reg [31:0] _RAND_26;
  reg  outputMemBlock_8;
  reg [31:0] _RAND_27;
  reg  outputMemBlock_9;
  reg [31:0] _RAND_28;
  reg  outputMemBlock_10;
  reg [31:0] _RAND_29;
  reg  outputMemBlock_11;
  reg [31:0] _RAND_30;
  reg  outputMemBlock_12;
  reg [31:0] _RAND_31;
  reg  outputMemBlock_13;
  reg [31:0] _RAND_32;
  reg  outputMemBlock_14;
  reg [31:0] _RAND_33;
  reg  outputMemBlock_15;
  reg [31:0] _RAND_34;
  reg [9:0] outputBits;
  reg [31:0] _RAND_35;
  reg [4:0] outputPieceBits;
  reg [31:0] _RAND_36;
  wire  inputBram_clock;
  wire [4:0] inputBram_io_a_addr;
  wire [15:0] inputBram_io_a_din;
  wire  inputBram_io_a_wr;
  wire [4:0] inputBram_io_b_addr;
  wire [15:0] inputBram_io_b_dout;
  reg [4:0] inputReadAddr;
  reg [31:0] _RAND_37;
  reg  inputPieceRead;
  reg [31:0] _RAND_38;
  wire  outputBram_clock;
  wire [4:0] outputBram_io_a_addr;
  wire [15:0] outputBram_io_a_din;
  wire  outputBram_io_a_wr;
  wire [4:0] outputBram_io_b_addr;
  wire [15:0] outputBram_io_b_dout;
  reg [4:0] outputWriteAddr;
  reg [31:0] _RAND_39;
  reg [4:0] outputReadAddr;
  reg [31:0] _RAND_40;
  wire  _T_75;
  wire  _T_76;
  wire  _GEN_0;
  wire [9:0] _GEN_1;
  wire  _T_79;
  wire  _T_80;
  wire  _GEN_2;
  wire  _T_84;
  wire  _T_85;
  wire  _T_89;
  wire  _T_90;
  wire  _T_92;
  wire  _T_96;
  wire [9:0] _T_98;
  wire [5:0] _T_100;
  wire [4:0] _T_101;
  wire  _T_102;
  wire  _T_103;
  wire  _T_104;
  wire  _T_105;
  wire  _T_106;
  wire  _T_107;
  wire  _T_108;
  wire  _T_109;
  wire  _T_110;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  _T_114;
  wire  _T_115;
  wire  _T_116;
  wire  _T_117;
  wire [9:0] _GEN_4;
  wire [4:0] _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [9:0] _GEN_23;
  wire [4:0] _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  inputAdvance;
  wire  _T_120;
  wire  _T_122;
  wire  _T_124;
  wire  _T_125;
  wire  _T_129;
  wire  _T_130;
  wire [5:0] _T_132;
  wire [5:0] _T_133;
  wire [4:0] _T_134;
  wire [10:0] _T_136;
  wire [10:0] _T_137;
  wire [9:0] _T_138;
  wire [9:0] _GEN_41;
  wire [9:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  nextBitValid;
  wire  nextBit;
  wire [5:0] _T_142;
  wire [4:0] _T_143;
  wire [10:0] _T_145;
  wire [9:0] _T_146;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire [4:0] _GEN_74;
  wire [9:0] _GEN_75;
  wire  _T_148;
  wire  _T_151;
  wire  _T_153;
  wire  _T_154;
  wire  _T_155;
  wire [1:0] _T_156;
  wire [1:0] _T_157;
  wire [3:0] _T_158;
  wire [1:0] _T_159;
  wire [1:0] _T_160;
  wire [3:0] _T_161;
  wire [7:0] _T_162;
  wire [1:0] _T_163;
  wire [1:0] _T_164;
  wire [3:0] _T_165;
  wire [1:0] _T_166;
  wire [1:0] _T_167;
  wire [3:0] _T_168;
  wire [7:0] _T_169;
  wire [15:0] _T_170;
  wire [5:0] _T_175;
  wire [4:0] _T_176;
  wire [4:0] _GEN_76;
  wire [4:0] _GEN_77;
  reg  outputReadingStarted;
  reg [31:0] _RAND_41;
  wire  _T_181;
  wire  _T_188;
  wire  _T_189;
  wire  _T_190;
  wire  _T_191;
  wire  _GEN_78;
  wire  _T_193;
  wire  _T_195;
  wire  _T_196;
  wire [5:0] _T_198;
  wire [4:0] _T_199;
  wire [4:0] _GEN_79;
  wire  _T_203;
  wire  _T_204;
  wire  _T_214;
  wire  _T_219;
  wire  _T_220;
  wire [9:0] _GEN_80;
  wire [4:0] _GEN_81;
  wire  _GEN_82;
  wire [4:0] _GEN_83;
  wire [4:0] _GEN_84;
  DualPortBRAM inputBram (
    .clock(inputBram_clock),
    .io_a_addr(inputBram_io_a_addr),
    .io_a_din(inputBram_io_a_din),
    .io_a_wr(inputBram_io_a_wr),
    .io_b_addr(inputBram_io_b_addr),
    .io_b_dout(inputBram_io_b_dout)
  );
  DualPortBRAM outputBram (
    .clock(outputBram_clock),
    .io_a_addr(outputBram_io_a_addr),
    .io_a_din(outputBram_io_a_din),
    .io_a_wr(outputBram_io_a_wr),
    .io_b_addr(outputBram_io_b_addr),
    .io_b_dout(outputBram_io_b_dout)
  );
  assign _T_75 = io_inputMemIdx == 5'h1f;
  assign _T_76 = io_inputMemBlockValid & _T_75;
  assign _GEN_0 = _T_76 ? 1'h1 : inputBlockLoaded;
  assign _GEN_1 = _T_76 ? io_inputBits : inputBitsRemaining;
  assign _T_79 = inputBitsRemaining == 10'h0;
  assign _T_80 = inputBlockLoaded & _T_79;
  assign _GEN_2 = _T_80 ? 1'h0 : _GEN_0;
  assign _T_84 = inputPieceBitsRemaining == 5'h0;
  assign _T_85 = inputBlockLoaded & _T_84;
  assign _T_89 = _T_79 == 1'h0;
  assign _T_90 = _T_85 & _T_89;
  assign _T_92 = inputPieceRead == 1'h0;
  assign _T_96 = inputBitsRemaining < 10'h10;
  assign _T_98 = _T_96 ? inputBitsRemaining : 10'h10;
  assign _T_100 = inputReadAddr + 5'h1;
  assign _T_101 = _T_100[4:0];
  assign _T_102 = inputBram_io_b_dout[0];
  assign _T_103 = inputBram_io_b_dout[1];
  assign _T_104 = inputBram_io_b_dout[2];
  assign _T_105 = inputBram_io_b_dout[3];
  assign _T_106 = inputBram_io_b_dout[4];
  assign _T_107 = inputBram_io_b_dout[5];
  assign _T_108 = inputBram_io_b_dout[6];
  assign _T_109 = inputBram_io_b_dout[7];
  assign _T_110 = inputBram_io_b_dout[8];
  assign _T_111 = inputBram_io_b_dout[9];
  assign _T_112 = inputBram_io_b_dout[10];
  assign _T_113 = inputBram_io_b_dout[11];
  assign _T_114 = inputBram_io_b_dout[12];
  assign _T_115 = inputBram_io_b_dout[13];
  assign _T_116 = inputBram_io_b_dout[14];
  assign _T_117 = inputBram_io_b_dout[15];
  assign _GEN_4 = _T_92 ? {{5'd0}, inputPieceBitsRemaining} : _T_98;
  assign _GEN_5 = _T_92 ? inputReadAddr : _T_101;
  assign _GEN_6 = _T_92 ? inputMemBlock_0 : _T_102;
  assign _GEN_7 = _T_92 ? inputMemBlock_1 : _T_103;
  assign _GEN_8 = _T_92 ? inputMemBlock_2 : _T_104;
  assign _GEN_9 = _T_92 ? inputMemBlock_3 : _T_105;
  assign _GEN_10 = _T_92 ? inputMemBlock_4 : _T_106;
  assign _GEN_11 = _T_92 ? inputMemBlock_5 : _T_107;
  assign _GEN_12 = _T_92 ? inputMemBlock_6 : _T_108;
  assign _GEN_13 = _T_92 ? inputMemBlock_7 : _T_109;
  assign _GEN_14 = _T_92 ? inputMemBlock_8 : _T_110;
  assign _GEN_15 = _T_92 ? inputMemBlock_9 : _T_111;
  assign _GEN_16 = _T_92 ? inputMemBlock_10 : _T_112;
  assign _GEN_17 = _T_92 ? inputMemBlock_11 : _T_113;
  assign _GEN_18 = _T_92 ? inputMemBlock_12 : _T_114;
  assign _GEN_19 = _T_92 ? inputMemBlock_13 : _T_115;
  assign _GEN_20 = _T_92 ? inputMemBlock_14 : _T_116;
  assign _GEN_21 = _T_92 ? inputMemBlock_15 : _T_117;
  assign _GEN_22 = _T_90 ? _T_92 : inputPieceRead;
  assign _GEN_23 = _T_90 ? _GEN_4 : {{5'd0}, inputPieceBitsRemaining};
  assign _GEN_24 = _T_90 ? _GEN_5 : inputReadAddr;
  assign _GEN_25 = _T_90 ? _GEN_6 : inputMemBlock_0;
  assign _GEN_26 = _T_90 ? _GEN_7 : inputMemBlock_1;
  assign _GEN_27 = _T_90 ? _GEN_8 : inputMemBlock_2;
  assign _GEN_28 = _T_90 ? _GEN_9 : inputMemBlock_3;
  assign _GEN_29 = _T_90 ? _GEN_10 : inputMemBlock_4;
  assign _GEN_30 = _T_90 ? _GEN_11 : inputMemBlock_5;
  assign _GEN_31 = _T_90 ? _GEN_12 : inputMemBlock_6;
  assign _GEN_32 = _T_90 ? _GEN_13 : inputMemBlock_7;
  assign _GEN_33 = _T_90 ? _GEN_14 : inputMemBlock_8;
  assign _GEN_34 = _T_90 ? _GEN_15 : inputMemBlock_9;
  assign _GEN_35 = _T_90 ? _GEN_16 : inputMemBlock_10;
  assign _GEN_36 = _T_90 ? _GEN_17 : inputMemBlock_11;
  assign _GEN_37 = _T_90 ? _GEN_18 : inputMemBlock_12;
  assign _GEN_38 = _T_90 ? _GEN_19 : inputMemBlock_13;
  assign _GEN_39 = _T_90 ? _GEN_20 : inputMemBlock_14;
  assign _GEN_40 = _T_90 ? _GEN_21 : inputMemBlock_15;
  assign _T_120 = outputPieceBits != 5'h10;
  assign _T_122 = outputBits == 10'h200;
  assign _T_124 = _T_122 == 1'h0;
  assign _T_125 = _T_120 & _T_124;
  assign _T_129 = _T_84 == 1'h0;
  assign _T_130 = _T_125 & _T_129;
  assign _T_132 = inputPieceBitsRemaining - 5'h1;
  assign _T_133 = $unsigned(_T_132);
  assign _T_134 = _T_133[4:0];
  assign _T_136 = inputBitsRemaining - 10'h1;
  assign _T_137 = $unsigned(_T_136);
  assign _T_138 = _T_137[9:0];
  assign _GEN_41 = inputAdvance ? {{5'd0}, _T_134} : _GEN_23;
  assign _GEN_42 = inputAdvance ? _T_138 : _GEN_1;
  assign _GEN_43 = inputAdvance ? inputMemBlock_1 : _GEN_25;
  assign _GEN_44 = inputAdvance ? inputMemBlock_2 : _GEN_26;
  assign _GEN_45 = inputAdvance ? inputMemBlock_3 : _GEN_27;
  assign _GEN_46 = inputAdvance ? inputMemBlock_4 : _GEN_28;
  assign _GEN_47 = inputAdvance ? inputMemBlock_5 : _GEN_29;
  assign _GEN_48 = inputAdvance ? inputMemBlock_6 : _GEN_30;
  assign _GEN_49 = inputAdvance ? inputMemBlock_7 : _GEN_31;
  assign _GEN_50 = inputAdvance ? inputMemBlock_8 : _GEN_32;
  assign _GEN_51 = inputAdvance ? inputMemBlock_9 : _GEN_33;
  assign _GEN_52 = inputAdvance ? inputMemBlock_10 : _GEN_34;
  assign _GEN_53 = inputAdvance ? inputMemBlock_11 : _GEN_35;
  assign _GEN_54 = inputAdvance ? inputMemBlock_12 : _GEN_36;
  assign _GEN_55 = inputAdvance ? inputMemBlock_13 : _GEN_37;
  assign _GEN_56 = inputAdvance ? inputMemBlock_14 : _GEN_38;
  assign _GEN_57 = inputAdvance ? inputMemBlock_15 : _GEN_39;
  assign _T_142 = outputPieceBits + 5'h1;
  assign _T_143 = _T_142[4:0];
  assign _T_145 = outputBits + 10'h1;
  assign _T_146 = _T_145[9:0];
  assign _GEN_58 = nextBitValid ? nextBit : outputMemBlock_15;
  assign _GEN_59 = nextBitValid ? outputMemBlock_1 : outputMemBlock_0;
  assign _GEN_60 = nextBitValid ? outputMemBlock_2 : outputMemBlock_1;
  assign _GEN_61 = nextBitValid ? outputMemBlock_3 : outputMemBlock_2;
  assign _GEN_62 = nextBitValid ? outputMemBlock_4 : outputMemBlock_3;
  assign _GEN_63 = nextBitValid ? outputMemBlock_5 : outputMemBlock_4;
  assign _GEN_64 = nextBitValid ? outputMemBlock_6 : outputMemBlock_5;
  assign _GEN_65 = nextBitValid ? outputMemBlock_7 : outputMemBlock_6;
  assign _GEN_66 = nextBitValid ? outputMemBlock_8 : outputMemBlock_7;
  assign _GEN_67 = nextBitValid ? outputMemBlock_9 : outputMemBlock_8;
  assign _GEN_68 = nextBitValid ? outputMemBlock_10 : outputMemBlock_9;
  assign _GEN_69 = nextBitValid ? outputMemBlock_11 : outputMemBlock_10;
  assign _GEN_70 = nextBitValid ? outputMemBlock_12 : outputMemBlock_11;
  assign _GEN_71 = nextBitValid ? outputMemBlock_13 : outputMemBlock_12;
  assign _GEN_72 = nextBitValid ? outputMemBlock_14 : outputMemBlock_13;
  assign _GEN_73 = nextBitValid ? outputMemBlock_15 : outputMemBlock_14;
  assign _GEN_74 = nextBitValid ? _T_143 : outputPieceBits;
  assign _GEN_75 = nextBitValid ? _T_146 : outputBits;
  assign _T_148 = outputPieceBits == 5'h10;
  assign _T_151 = io_inputFinished & _T_79;
  assign _T_153 = outputPieceBits > 5'h0;
  assign _T_154 = _T_151 & _T_153;
  assign _T_155 = _T_148 | _T_154;
  assign _T_156 = {outputMemBlock_1,outputMemBlock_0};
  assign _T_157 = {outputMemBlock_3,outputMemBlock_2};
  assign _T_158 = {_T_157,_T_156};
  assign _T_159 = {outputMemBlock_5,outputMemBlock_4};
  assign _T_160 = {outputMemBlock_7,outputMemBlock_6};
  assign _T_161 = {_T_160,_T_159};
  assign _T_162 = {_T_161,_T_158};
  assign _T_163 = {outputMemBlock_9,outputMemBlock_8};
  assign _T_164 = {outputMemBlock_11,outputMemBlock_10};
  assign _T_165 = {_T_164,_T_163};
  assign _T_166 = {outputMemBlock_13,outputMemBlock_12};
  assign _T_167 = {outputMemBlock_15,outputMemBlock_14};
  assign _T_168 = {_T_167,_T_166};
  assign _T_169 = {_T_168,_T_165};
  assign _T_170 = {_T_169,_T_162};
  assign _T_175 = outputWriteAddr + 5'h1;
  assign _T_176 = _T_175[4:0];
  assign _GEN_76 = _T_148 ? 5'h0 : _GEN_74;
  assign _GEN_77 = _T_148 ? _T_176 : outputWriteAddr;
  assign _T_181 = outputReadingStarted == 1'h0;
  assign _T_188 = outputBits > 10'h0;
  assign _T_189 = _T_151 & _T_188;
  assign _T_190 = _T_122 | _T_189;
  assign _T_191 = _T_181 & _T_190;
  assign _GEN_78 = _T_191 ? 1'h1 : outputReadingStarted;
  assign _T_193 = io_outputMemBlockReady & outputReadingStarted;
  assign _T_195 = outputReadAddr != 5'h1f;
  assign _T_196 = _T_193 & _T_195;
  assign _T_198 = outputReadAddr + 5'h1;
  assign _T_199 = _T_198[4:0];
  assign _GEN_79 = _T_196 ? _T_199 : outputReadAddr;
  assign _T_203 = io_inputFinished == 1'h0;
  assign _T_204 = _T_79 & _T_203;
  assign _T_214 = outputReadingStarted & _T_190;
  assign _T_219 = outputBits == 10'h0;
  assign _T_220 = _T_151 & _T_219;
  assign _GEN_80 = io_outputMemFlushed ? 10'h0 : _GEN_75;
  assign _GEN_81 = io_outputMemFlushed ? 5'h0 : _GEN_76;
  assign _GEN_82 = io_outputMemFlushed ? 1'h0 : _GEN_78;
  assign _GEN_83 = io_outputMemFlushed ? 5'h0 : _GEN_77;
  assign _GEN_84 = io_outputMemFlushed ? 5'h0 : _GEN_79;
  assign io_inputMemConsumed = _T_204;
  assign io_outputMemBlock = outputBram_io_b_dout;
  assign io_outputMemBlockValid = _T_214;
  assign io_outputBits = outputBits;
  assign io_outputFinished = _T_220;
  assign inputBram_io_a_addr = io_inputMemIdx;
  assign inputBram_io_a_din = io_inputMemBlock;
  assign inputBram_io_a_wr = io_inputMemBlockValid;
  assign inputBram_io_b_addr = inputReadAddr;
  assign inputBram_clock = clock;
  assign outputBram_io_a_addr = outputWriteAddr;
  assign outputBram_io_a_din = _T_170;
  assign outputBram_io_a_wr = _T_155;
  assign outputBram_io_b_addr = outputReadAddr;
  assign outputBram_clock = clock;
  assign inputAdvance = _T_130;
  assign nextBitValid = inputAdvance;
  assign nextBit = inputMemBlock_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  inputMemBlock_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  inputMemBlock_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputMemBlock_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  inputMemBlock_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  inputMemBlock_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  inputMemBlock_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  inputMemBlock_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemBlock_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBlock_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  inputMemBlock_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputMemBlock_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  inputMemBlock_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  inputMemBlock_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  inputMemBlock_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  inputMemBlock_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  inputMemBlock_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  inputPieceBitsRemaining = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  inputBitsRemaining = _RAND_17[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  inputBlockLoaded = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  outputMemBlock_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  outputMemBlock_1 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  outputMemBlock_2 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  outputMemBlock_3 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  outputMemBlock_4 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  outputMemBlock_5 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  outputMemBlock_6 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  outputMemBlock_7 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  outputMemBlock_8 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  outputMemBlock_9 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  outputMemBlock_10 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  outputMemBlock_11 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  outputMemBlock_12 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  outputMemBlock_13 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  outputMemBlock_14 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  outputMemBlock_15 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  outputBits = _RAND_35[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  outputPieceBits = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  inputReadAddr = _RAND_37[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  inputPieceRead = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  outputWriteAddr = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  outputReadAddr = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  outputReadingStarted = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (inputAdvance) begin
      inputMemBlock_0 <= inputMemBlock_1;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_0 <= _T_102;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_1 <= inputMemBlock_2;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_1 <= _T_103;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_2 <= inputMemBlock_3;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_2 <= _T_104;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_3 <= inputMemBlock_4;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_3 <= _T_105;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_4 <= inputMemBlock_5;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_4 <= _T_106;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_5 <= inputMemBlock_6;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_5 <= _T_107;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_6 <= inputMemBlock_7;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_6 <= _T_108;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_7 <= inputMemBlock_8;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_7 <= _T_109;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_8 <= inputMemBlock_9;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_8 <= _T_110;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_9 <= inputMemBlock_10;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_9 <= _T_111;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_10 <= inputMemBlock_11;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_10 <= _T_112;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_11 <= inputMemBlock_12;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_11 <= _T_113;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_12 <= inputMemBlock_13;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_12 <= _T_114;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_13 <= inputMemBlock_14;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_13 <= _T_115;
        end
      end
    end
    if (inputAdvance) begin
      inputMemBlock_14 <= inputMemBlock_15;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputMemBlock_14 <= _T_116;
        end
      end
    end
    if (_T_90) begin
      if (!(_T_92)) begin
        inputMemBlock_15 <= _T_117;
      end
    end
    if (reset) begin
      inputPieceBitsRemaining <= 5'h0;
    end else begin
      inputPieceBitsRemaining <= _GEN_41[4:0];
    end
    if (reset) begin
      inputBitsRemaining <= 10'h0;
    end else begin
      if (inputAdvance) begin
        inputBitsRemaining <= _T_138;
      end else begin
        if (_T_76) begin
          inputBitsRemaining <= io_inputBits;
        end
      end
    end
    if (reset) begin
      inputBlockLoaded <= 1'h0;
    end else begin
      if (_T_80) begin
        inputBlockLoaded <= 1'h0;
      end else begin
        if (_T_76) begin
          inputBlockLoaded <= 1'h1;
        end
      end
    end
    if (nextBitValid) begin
      outputMemBlock_0 <= outputMemBlock_1;
    end
    if (nextBitValid) begin
      outputMemBlock_1 <= outputMemBlock_2;
    end
    if (nextBitValid) begin
      outputMemBlock_2 <= outputMemBlock_3;
    end
    if (nextBitValid) begin
      outputMemBlock_3 <= outputMemBlock_4;
    end
    if (nextBitValid) begin
      outputMemBlock_4 <= outputMemBlock_5;
    end
    if (nextBitValid) begin
      outputMemBlock_5 <= outputMemBlock_6;
    end
    if (nextBitValid) begin
      outputMemBlock_6 <= outputMemBlock_7;
    end
    if (nextBitValid) begin
      outputMemBlock_7 <= outputMemBlock_8;
    end
    if (nextBitValid) begin
      outputMemBlock_8 <= outputMemBlock_9;
    end
    if (nextBitValid) begin
      outputMemBlock_9 <= outputMemBlock_10;
    end
    if (nextBitValid) begin
      outputMemBlock_10 <= outputMemBlock_11;
    end
    if (nextBitValid) begin
      outputMemBlock_11 <= outputMemBlock_12;
    end
    if (nextBitValid) begin
      outputMemBlock_12 <= outputMemBlock_13;
    end
    if (nextBitValid) begin
      outputMemBlock_13 <= outputMemBlock_14;
    end
    if (nextBitValid) begin
      outputMemBlock_14 <= outputMemBlock_15;
    end
    if (nextBitValid) begin
      outputMemBlock_15 <= nextBit;
    end
    if (reset) begin
      outputBits <= 10'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputBits <= 10'h0;
      end else begin
        if (nextBitValid) begin
          outputBits <= _T_146;
        end
      end
    end
    if (reset) begin
      outputPieceBits <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputPieceBits <= 5'h0;
      end else begin
        if (_T_148) begin
          outputPieceBits <= 5'h0;
        end else begin
          if (nextBitValid) begin
            outputPieceBits <= _T_143;
          end
        end
      end
    end
    if (reset) begin
      inputReadAddr <= 5'h0;
    end else begin
      if (_T_90) begin
        if (!(_T_92)) begin
          inputReadAddr <= _T_101;
        end
      end
    end
    if (reset) begin
      inputPieceRead <= 1'h0;
    end else begin
      if (_T_90) begin
        inputPieceRead <= _T_92;
      end
    end
    if (reset) begin
      outputWriteAddr <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputWriteAddr <= 5'h0;
      end else begin
        if (_T_148) begin
          outputWriteAddr <= _T_176;
        end
      end
    end
    if (reset) begin
      outputReadAddr <= 5'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputReadAddr <= 5'h0;
      end else begin
        if (_T_196) begin
          outputReadAddr <= _T_199;
        end
      end
    end
    if (reset) begin
      outputReadingStarted <= 1'h0;
    end else begin
      if (io_outputMemFlushed) begin
        outputReadingStarted <= 1'h0;
      end else begin
        if (_T_191) begin
          outputReadingStarted <= 1'h1;
        end
      end
    end
  end
endmodule
module StreamingCore(
  input         clock,
  input         reset,
  output [31:0] io_inputMemAddr,
  input         io_inputMemAddrConsumed,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output        io_inputMemBlockReady,
  output [31:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [15:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output        io_inputAddrsIgnore,
  output        io_inputBlocksFinished,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [15:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [15:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [31:0] inputBitsRemaining;
  reg [31:0] _RAND_2;
  reg  coreInputFinished;
  reg [31:0] _RAND_3;
  reg [31:0] outputBits;
  reg [31:0] _RAND_4;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_5;
  reg  outputLengthCommitted;
  reg [31:0] _RAND_6;
  reg [31:0] inputMemAddr;
  reg [31:0] _RAND_7;
  reg [31:0] inputMemBound;
  reg [31:0] _RAND_8;
  reg [31:0] outputMemAddr;
  reg [31:0] _RAND_9;
  reg [31:0] outputLenAddr;
  reg [31:0] _RAND_10;
  wire  _T_40;
  wire  _T_41;
  wire  _T_44;
  reg  initAddressAcked;
  reg [31:0] _RAND_11;
  wire  _GEN_0;
  wire  _T_48;
  wire [32:0] _T_50;
  wire [31:0] _T_51;
  wire [31:0] _GEN_1;
  wire  _T_52;
  wire  _T_53;
  wire  _T_54;
  wire  _T_55;
  wire  _T_56;
  wire  _T_58;
  wire  _T_60;
  wire  _T_61;
  wire  _T_62;
  wire  _T_63;
  wire  _T_65;
  wire [31:0] _T_67;
  wire  _T_69;
  wire [15:0] _T_70;
  wire [31:0] _T_71;
  wire [31:0] _GEN_2;
  wire  _T_73;
  wire [15:0] _T_74;
  wire [31:0] _T_75;
  wire [31:0] _GEN_3;
  wire  _T_77;
  wire [15:0] _T_78;
  wire [31:0] _T_79;
  wire [22:0] _T_80;
  wire [28:0] _T_82;
  wire [31:0] _GEN_44;
  wire [32:0] _T_83;
  wire [31:0] _T_84;
  wire [8:0] _T_85;
  wire  _T_87;
  wire [6:0] _T_90;
  wire [31:0] _GEN_45;
  wire [32:0] _T_91;
  wire [31:0] _T_92;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire  _T_94;
  wire [15:0] _T_95;
  wire [31:0] _T_96;
  wire [22:0] _T_97;
  wire [28:0] _T_99;
  wire [31:0] _GEN_46;
  wire [32:0] _T_100;
  wire [31:0] _T_101;
  wire [8:0] _T_102;
  wire  _T_104;
  wire [6:0] _T_107;
  wire [31:0] _GEN_47;
  wire [32:0] _T_108;
  wire [31:0] _T_109;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire  _T_111;
  wire [15:0] _T_112;
  wire [31:0] _T_113;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire  _T_115;
  wire [15:0] _T_116;
  wire [31:0] _T_117;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire  _T_119;
  wire [32:0] _T_123;
  wire [31:0] _T_124;
  wire  _GEN_12;
  wire  _GEN_13;
  wire [31:0] _GEN_14;
  wire [32:0] _T_130;
  wire [32:0] _T_131;
  wire [31:0] _T_132;
  wire [31:0] _T_134;
  wire [31:0] _GEN_15;
  wire [31:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [31:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [31:0] _GEN_23;
  wire [31:0] _GEN_24;
  wire [31:0] _GEN_25;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _T_139;
  wire  _GEN_30;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_12;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_13;
  wire  _GEN_31;
  wire [31:0] _T_146;
  wire  _T_148;
  wire  _T_150;
  wire  _T_151;
  wire  _T_152;
  wire  _T_153;
  wire  _T_154;
  wire  _GEN_32;
  wire  _T_160;
  wire [4:0] _GEN_33;
  wire [5:0] _T_163;
  wire [4:0] _T_164;
  wire [4:0] _GEN_34;
  wire [4:0] _GEN_35;
  wire [15:0] outputBitsBlock;
  wire  _T_167;
  wire [15:0] _T_168;
  wire  _T_170;
  wire [15:0] _T_171;
  wire [15:0] _T_173;
  wire [15:0] _T_174;
  wire [15:0] _T_175;
  wire  _T_176;
  wire  _T_180;
  wire [31:0] _GEN_48;
  wire [32:0] _T_184;
  wire [31:0] _T_185;
  wire  _GEN_36;
  wire [31:0] _GEN_37;
  wire [31:0] _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign _T_40 = io_inputAddrsIgnore == 1'h0;
  assign _T_41 = io_inputMemAddrConsumed & _T_40;
  assign _T_44 = reset == 1'h0;
  assign _GEN_0 = io_inputMemAddrConsumed ? 1'h1 : initAddressAcked;
  assign _T_48 = io_inputMemAddrConsumed & initDone;
  assign _T_50 = inputMemAddr + 32'h40;
  assign _T_51 = _T_50[31:0];
  assign _GEN_1 = _T_48 ? _T_51 : inputMemAddr;
  assign _T_52 = isInit & initAddressAcked;
  assign _T_53 = inputMemAddr == inputMemBound;
  assign _T_54 = initDone & _T_53;
  assign _T_55 = _T_52 | _T_54;
  assign _T_56 = initDone & core_io_inputMemConsumed;
  assign _T_58 = inputBitsRemaining == 32'h0;
  assign _T_60 = _T_58 == 1'h0;
  assign _T_61 = _T_56 & _T_60;
  assign _T_62 = isInit | _T_61;
  assign _T_63 = io_inputMemBlockValid & initDone;
  assign _T_65 = inputBitsRemaining > 32'h200;
  assign _T_67 = _T_65 ? 32'h200 : inputBitsRemaining;
  assign _T_69 = io_inputMemIdx == 5'h0;
  assign _T_70 = inputMemAddr[31:16];
  assign _T_71 = {_T_70,io_inputMemBlock};
  assign _GEN_2 = _T_69 ? _T_71 : _GEN_1;
  assign _T_73 = io_inputMemIdx == 5'h1;
  assign _T_74 = inputMemAddr[15:0];
  assign _T_75 = {io_inputMemBlock,_T_74};
  assign _GEN_3 = _T_73 ? _T_75 : _GEN_2;
  assign _T_77 = io_inputMemIdx == 5'h4;
  assign _T_78 = inputBitsRemaining[31:16];
  assign _T_79 = {_T_78,io_inputMemBlock};
  assign _T_80 = _T_79[31:9];
  assign _T_82 = {_T_80,6'h0};
  assign _GEN_44 = {{3'd0}, _T_82};
  assign _T_83 = inputMemAddr + _GEN_44;
  assign _T_84 = _T_83[31:0];
  assign _T_85 = _T_79[8:0];
  assign _T_87 = _T_85 != 9'h0;
  assign _T_90 = _T_87 ? 7'h40 : 7'h0;
  assign _GEN_45 = {{25'd0}, _T_90};
  assign _T_91 = _T_84 + _GEN_45;
  assign _T_92 = _T_91[31:0];
  assign _GEN_4 = _T_77 ? _T_79 : inputBitsRemaining;
  assign _GEN_5 = _T_77 ? _T_92 : inputMemBound;
  assign _T_94 = io_inputMemIdx == 5'h5;
  assign _T_95 = inputBitsRemaining[15:0];
  assign _T_96 = {io_inputMemBlock,_T_95};
  assign _T_97 = _T_96[31:9];
  assign _T_99 = {_T_97,6'h0};
  assign _GEN_46 = {{3'd0}, _T_99};
  assign _T_100 = inputMemAddr + _GEN_46;
  assign _T_101 = _T_100[31:0];
  assign _T_102 = _T_96[8:0];
  assign _T_104 = _T_102 != 9'h0;
  assign _T_107 = _T_104 ? 7'h40 : 7'h0;
  assign _GEN_47 = {{25'd0}, _T_107};
  assign _T_108 = _T_101 + _GEN_47;
  assign _T_109 = _T_108[31:0];
  assign _GEN_6 = _T_94 ? _T_96 : _GEN_4;
  assign _GEN_7 = _T_94 ? _T_109 : _GEN_5;
  assign _T_111 = io_inputMemIdx == 5'h8;
  assign _T_112 = outputMemAddr[31:16];
  assign _T_113 = {_T_112,io_inputMemBlock};
  assign _GEN_8 = _T_111 ? _T_113 : outputMemAddr;
  assign _GEN_9 = _T_111 ? _T_113 : outputLenAddr;
  assign _T_115 = io_inputMemIdx == 5'h9;
  assign _T_116 = outputMemAddr[15:0];
  assign _T_117 = {io_inputMemBlock,_T_116};
  assign _GEN_10 = _T_115 ? _T_117 : _GEN_8;
  assign _GEN_11 = _T_115 ? _T_117 : _GEN_9;
  assign _T_119 = io_inputMemIdx == 5'h1f;
  assign _T_123 = outputMemAddr + 32'h40;
  assign _T_124 = _T_123[31:0];
  assign _GEN_12 = _T_119 ? 1'h0 : isInit;
  assign _GEN_13 = _T_119 ? 1'h1 : initDone;
  assign _GEN_14 = _T_119 ? _T_124 : _GEN_10;
  assign _T_130 = inputBitsRemaining - 32'h200;
  assign _T_131 = $unsigned(_T_130);
  assign _T_132 = _T_131[31:0];
  assign _T_134 = _T_65 ? _T_132 : 32'h0;
  assign _GEN_15 = _T_119 ? _T_134 : inputBitsRemaining;
  assign _GEN_16 = isInit ? _GEN_3 : _GEN_1;
  assign _GEN_17 = isInit ? _GEN_6 : _GEN_15;
  assign _GEN_18 = isInit ? _GEN_7 : inputMemBound;
  assign _GEN_19 = isInit ? _GEN_14 : outputMemAddr;
  assign _GEN_20 = isInit ? _GEN_11 : outputLenAddr;
  assign _GEN_21 = isInit ? _GEN_12 : isInit;
  assign _GEN_22 = isInit ? _GEN_13 : initDone;
  assign _GEN_23 = io_inputMemBlockValid ? _GEN_16 : _GEN_1;
  assign _GEN_24 = io_inputMemBlockValid ? _GEN_17 : inputBitsRemaining;
  assign _GEN_25 = io_inputMemBlockValid ? _GEN_18 : inputMemBound;
  assign _GEN_26 = io_inputMemBlockValid ? _GEN_19 : outputMemAddr;
  assign _GEN_27 = io_inputMemBlockValid ? _GEN_20 : outputLenAddr;
  assign _GEN_28 = io_inputMemBlockValid ? _GEN_21 : isInit;
  assign _GEN_29 = io_inputMemBlockValid ? _GEN_22 : initDone;
  assign _T_139 = core_io_inputMemConsumed & _T_58;
  assign _GEN_30 = _T_139 ? 1'h1 : coreInputFinished;
  assign _GEN_31 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_146 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_148 = outputAddressAccepted == 1'h0;
  assign _T_150 = outputLengthCommitted == 1'h0;
  assign _T_151 = core_io_outputFinished & _T_150;
  assign _T_152 = core_io_outputMemBlockValid | _T_151;
  assign _T_153 = _T_148 & _T_152;
  assign _T_154 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_32 = _T_154 ? 1'h1 : outputAddressAccepted;
  assign _T_160 = outputBlockCounter == 5'h1f;
  assign _GEN_33 = io_outputMemBlockReady ? 5'h0 : outputBlockCounter;
  assign _T_163 = outputBlockCounter + 5'h1;
  assign _T_164 = _T_163[4:0];
  assign _GEN_34 = _T_160 ? _GEN_33 : _T_164;
  assign _GEN_35 = outputAddressAcceptedNext ? _GEN_34 : outputBlockCounter;
  assign _T_167 = outputBlockCounter == 5'h0;
  assign _T_168 = outputBits[15:0];
  assign _T_170 = outputBlockCounter == 5'h1;
  assign _T_171 = outputBits[31:16];
  assign _T_173 = _T_170 ? _T_171 : 16'h0;
  assign _T_174 = _T_167 ? _T_168 : _T_173;
  assign _T_175 = core_io_outputFinished ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_176 = outputAddressAcceptedNext & io_outputMemBlockReady;
  assign _T_180 = _T_176 & _T_160;
  assign _GEN_48 = {{22'd0}, core_io_outputBits};
  assign _T_184 = outputBits + _GEN_48;
  assign _T_185 = _T_184[31:0];
  assign _GEN_36 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _GEN_37 = core_io_outputFinished ? outputBits : _T_185;
  assign _GEN_38 = core_io_outputFinished ? _GEN_26 : _T_124;
  assign _GEN_39 = _T_180 ? 1'h0 : _GEN_32;
  assign _GEN_40 = _T_180 ? 1'h0 : _GEN_31;
  assign _GEN_41 = _T_180 ? _GEN_36 : outputLengthCommitted;
  assign _GEN_42 = _T_180 ? _GEN_37 : outputBits;
  assign _GEN_43 = _T_180 ? _GEN_38 : _GEN_26;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemBlockReady = _T_62;
  assign io_outputMemAddr = _T_146;
  assign io_outputMemAddrValid = _T_153;
  assign io_outputMemBlock = _T_175;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_inputAddrsIgnore = _T_55;
  assign io_inputBlocksFinished = _T_58;
  assign io_outputFinished = outputLengthCommitted;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_63;
  assign core_io_inputBits = _T_67[9:0];
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_io_outputMemFlushed = _T_176;
  assign core_clock = clock;
  assign core_reset = reset;
  assign outputBitsBlock = _T_174;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputBitsRemaining = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  coreInputFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  outputBits = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputBlockCounter = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputLengthCommitted = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemAddr = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBound = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  outputMemAddr = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  outputLenAddr = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  initAddressAcked = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  outputAddressAccepted = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  outputAddressAcceptedNext = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_119) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_119) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 32'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_94) begin
            inputBitsRemaining <= _T_96;
          end else begin
            if (_T_77) begin
              inputBitsRemaining <= _T_79;
            end
          end
        end else begin
          if (_T_119) begin
            if (_T_65) begin
              inputBitsRemaining <= _T_132;
            end else begin
              inputBitsRemaining <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_139) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 32'h0;
    end else begin
      if (_T_180) begin
        if (!(core_io_outputFinished)) begin
          outputBits <= _T_185;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_160) begin
          if (io_outputMemBlockReady) begin
            outputBlockCounter <= 5'h0;
          end
        end else begin
          outputBlockCounter <= _T_164;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_180) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 32'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_73) begin
            inputMemAddr <= _T_75;
          end else begin
            if (_T_69) begin
              inputMemAddr <= _T_71;
            end else begin
              if (_T_48) begin
                inputMemAddr <= _T_51;
              end
            end
          end
        end else begin
          if (_T_48) begin
            inputMemAddr <= _T_51;
          end
        end
      end else begin
        if (_T_48) begin
          inputMemAddr <= _T_51;
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_94) begin
          inputMemBound <= _T_109;
        end else begin
          if (_T_77) begin
            inputMemBound <= _T_92;
          end
        end
      end
    end
    if (_T_180) begin
      if (core_io_outputFinished) begin
        if (io_inputMemBlockValid) begin
          if (isInit) begin
            if (_T_119) begin
              outputMemAddr <= _T_124;
            end else begin
              if (_T_115) begin
                outputMemAddr <= _T_117;
              end else begin
                if (_T_111) begin
                  outputMemAddr <= _T_113;
                end
              end
            end
          end
        end
      end else begin
        outputMemAddr <= _T_124;
      end
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_119) begin
            outputMemAddr <= _T_124;
          end else begin
            if (_T_115) begin
              outputMemAddr <= _T_117;
            end else begin
              if (_T_111) begin
                outputMemAddr <= _T_113;
              end
            end
          end
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_115) begin
          outputLenAddr <= _T_117;
        end else begin
          if (_T_111) begin
            outputLenAddr <= _T_113;
          end
        end
      end
    end
    if (reset) begin
      initAddressAcked <= 1'h0;
    end else begin
      if (io_inputMemAddrConsumed) begin
        initAddressAcked <= 1'h1;
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_180) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_154) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_180) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41 & _T_44) begin
          $fwrite(32'h80000002,"input address 0x%h accepted for core 0\n",io_inputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_154 & _T_44) begin
          $fwrite(32'h80000002,"output address 0x%h accepted for core 0\n",io_outputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module StreamingCore_1(
  input         clock,
  input         reset,
  output [31:0] io_inputMemAddr,
  input         io_inputMemAddrConsumed,
  input  [15:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output        io_inputMemBlockReady,
  output [31:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [15:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output        io_inputAddrsIgnore,
  output        io_inputBlocksFinished,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [15:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [9:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [15:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [9:0] core_io_outputBits;
  wire  core_io_outputFinished;
  wire  core_io_outputMemFlushed;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [31:0] inputBitsRemaining;
  reg [31:0] _RAND_2;
  reg  coreInputFinished;
  reg [31:0] _RAND_3;
  reg [31:0] outputBits;
  reg [31:0] _RAND_4;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_5;
  reg  outputLengthCommitted;
  reg [31:0] _RAND_6;
  reg [31:0] inputMemAddr;
  reg [31:0] _RAND_7;
  reg [31:0] inputMemBound;
  reg [31:0] _RAND_8;
  reg [31:0] outputMemAddr;
  reg [31:0] _RAND_9;
  reg [31:0] outputLenAddr;
  reg [31:0] _RAND_10;
  wire  _T_40;
  wire  _T_41;
  wire  _T_44;
  reg  initAddressAcked;
  reg [31:0] _RAND_11;
  wire  _GEN_0;
  wire  _T_48;
  wire [32:0] _T_50;
  wire [31:0] _T_51;
  wire [31:0] _GEN_1;
  wire  _T_52;
  wire  _T_53;
  wire  _T_54;
  wire  _T_55;
  wire  _T_56;
  wire  _T_58;
  wire  _T_60;
  wire  _T_61;
  wire  _T_62;
  wire  _T_63;
  wire  _T_65;
  wire [31:0] _T_67;
  wire  _T_69;
  wire [15:0] _T_70;
  wire [31:0] _T_71;
  wire [31:0] _GEN_2;
  wire  _T_73;
  wire [15:0] _T_74;
  wire [31:0] _T_75;
  wire [31:0] _GEN_3;
  wire  _T_77;
  wire [15:0] _T_78;
  wire [31:0] _T_79;
  wire [22:0] _T_80;
  wire [28:0] _T_82;
  wire [31:0] _GEN_44;
  wire [32:0] _T_83;
  wire [31:0] _T_84;
  wire [8:0] _T_85;
  wire  _T_87;
  wire [6:0] _T_90;
  wire [31:0] _GEN_45;
  wire [32:0] _T_91;
  wire [31:0] _T_92;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire  _T_94;
  wire [15:0] _T_95;
  wire [31:0] _T_96;
  wire [22:0] _T_97;
  wire [28:0] _T_99;
  wire [31:0] _GEN_46;
  wire [32:0] _T_100;
  wire [31:0] _T_101;
  wire [8:0] _T_102;
  wire  _T_104;
  wire [6:0] _T_107;
  wire [31:0] _GEN_47;
  wire [32:0] _T_108;
  wire [31:0] _T_109;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire  _T_111;
  wire [15:0] _T_112;
  wire [31:0] _T_113;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire  _T_115;
  wire [15:0] _T_116;
  wire [31:0] _T_117;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire  _T_119;
  wire [32:0] _T_123;
  wire [31:0] _T_124;
  wire  _GEN_12;
  wire  _GEN_13;
  wire [31:0] _GEN_14;
  wire [32:0] _T_130;
  wire [32:0] _T_131;
  wire [31:0] _T_132;
  wire [31:0] _T_134;
  wire [31:0] _GEN_15;
  wire [31:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [31:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire [31:0] _GEN_23;
  wire [31:0] _GEN_24;
  wire [31:0] _GEN_25;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _T_139;
  wire  _GEN_30;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_12;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_13;
  wire  _GEN_31;
  wire [31:0] _T_146;
  wire  _T_148;
  wire  _T_150;
  wire  _T_151;
  wire  _T_152;
  wire  _T_153;
  wire  _T_154;
  wire  _GEN_32;
  wire  _T_160;
  wire [4:0] _GEN_33;
  wire [5:0] _T_163;
  wire [4:0] _T_164;
  wire [4:0] _GEN_34;
  wire [4:0] _GEN_35;
  wire [15:0] outputBitsBlock;
  wire  _T_167;
  wire [15:0] _T_168;
  wire  _T_170;
  wire [15:0] _T_171;
  wire [15:0] _T_173;
  wire [15:0] _T_174;
  wire [15:0] _T_175;
  wire  _T_176;
  wire  _T_180;
  wire [31:0] _GEN_48;
  wire [32:0] _T_184;
  wire [31:0] _T_185;
  wire  _GEN_36;
  wire [31:0] _GEN_37;
  wire [31:0] _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  PassThrough core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished),
    .io_outputMemFlushed(core_io_outputMemFlushed)
  );
  assign _T_40 = io_inputAddrsIgnore == 1'h0;
  assign _T_41 = io_inputMemAddrConsumed & _T_40;
  assign _T_44 = reset == 1'h0;
  assign _GEN_0 = io_inputMemAddrConsumed ? 1'h1 : initAddressAcked;
  assign _T_48 = io_inputMemAddrConsumed & initDone;
  assign _T_50 = inputMemAddr + 32'h40;
  assign _T_51 = _T_50[31:0];
  assign _GEN_1 = _T_48 ? _T_51 : inputMemAddr;
  assign _T_52 = isInit & initAddressAcked;
  assign _T_53 = inputMemAddr == inputMemBound;
  assign _T_54 = initDone & _T_53;
  assign _T_55 = _T_52 | _T_54;
  assign _T_56 = initDone & core_io_inputMemConsumed;
  assign _T_58 = inputBitsRemaining == 32'h0;
  assign _T_60 = _T_58 == 1'h0;
  assign _T_61 = _T_56 & _T_60;
  assign _T_62 = isInit | _T_61;
  assign _T_63 = io_inputMemBlockValid & initDone;
  assign _T_65 = inputBitsRemaining > 32'h200;
  assign _T_67 = _T_65 ? 32'h200 : inputBitsRemaining;
  assign _T_69 = io_inputMemIdx == 5'h0;
  assign _T_70 = inputMemAddr[31:16];
  assign _T_71 = {_T_70,io_inputMemBlock};
  assign _GEN_2 = _T_69 ? _T_71 : _GEN_1;
  assign _T_73 = io_inputMemIdx == 5'h1;
  assign _T_74 = inputMemAddr[15:0];
  assign _T_75 = {io_inputMemBlock,_T_74};
  assign _GEN_3 = _T_73 ? _T_75 : _GEN_2;
  assign _T_77 = io_inputMemIdx == 5'h4;
  assign _T_78 = inputBitsRemaining[31:16];
  assign _T_79 = {_T_78,io_inputMemBlock};
  assign _T_80 = _T_79[31:9];
  assign _T_82 = {_T_80,6'h0};
  assign _GEN_44 = {{3'd0}, _T_82};
  assign _T_83 = inputMemAddr + _GEN_44;
  assign _T_84 = _T_83[31:0];
  assign _T_85 = _T_79[8:0];
  assign _T_87 = _T_85 != 9'h0;
  assign _T_90 = _T_87 ? 7'h40 : 7'h0;
  assign _GEN_45 = {{25'd0}, _T_90};
  assign _T_91 = _T_84 + _GEN_45;
  assign _T_92 = _T_91[31:0];
  assign _GEN_4 = _T_77 ? _T_79 : inputBitsRemaining;
  assign _GEN_5 = _T_77 ? _T_92 : inputMemBound;
  assign _T_94 = io_inputMemIdx == 5'h5;
  assign _T_95 = inputBitsRemaining[15:0];
  assign _T_96 = {io_inputMemBlock,_T_95};
  assign _T_97 = _T_96[31:9];
  assign _T_99 = {_T_97,6'h0};
  assign _GEN_46 = {{3'd0}, _T_99};
  assign _T_100 = inputMemAddr + _GEN_46;
  assign _T_101 = _T_100[31:0];
  assign _T_102 = _T_96[8:0];
  assign _T_104 = _T_102 != 9'h0;
  assign _T_107 = _T_104 ? 7'h40 : 7'h0;
  assign _GEN_47 = {{25'd0}, _T_107};
  assign _T_108 = _T_101 + _GEN_47;
  assign _T_109 = _T_108[31:0];
  assign _GEN_6 = _T_94 ? _T_96 : _GEN_4;
  assign _GEN_7 = _T_94 ? _T_109 : _GEN_5;
  assign _T_111 = io_inputMemIdx == 5'h8;
  assign _T_112 = outputMemAddr[31:16];
  assign _T_113 = {_T_112,io_inputMemBlock};
  assign _GEN_8 = _T_111 ? _T_113 : outputMemAddr;
  assign _GEN_9 = _T_111 ? _T_113 : outputLenAddr;
  assign _T_115 = io_inputMemIdx == 5'h9;
  assign _T_116 = outputMemAddr[15:0];
  assign _T_117 = {io_inputMemBlock,_T_116};
  assign _GEN_10 = _T_115 ? _T_117 : _GEN_8;
  assign _GEN_11 = _T_115 ? _T_117 : _GEN_9;
  assign _T_119 = io_inputMemIdx == 5'h1f;
  assign _T_123 = outputMemAddr + 32'h40;
  assign _T_124 = _T_123[31:0];
  assign _GEN_12 = _T_119 ? 1'h0 : isInit;
  assign _GEN_13 = _T_119 ? 1'h1 : initDone;
  assign _GEN_14 = _T_119 ? _T_124 : _GEN_10;
  assign _T_130 = inputBitsRemaining - 32'h200;
  assign _T_131 = $unsigned(_T_130);
  assign _T_132 = _T_131[31:0];
  assign _T_134 = _T_65 ? _T_132 : 32'h0;
  assign _GEN_15 = _T_119 ? _T_134 : inputBitsRemaining;
  assign _GEN_16 = isInit ? _GEN_3 : _GEN_1;
  assign _GEN_17 = isInit ? _GEN_6 : _GEN_15;
  assign _GEN_18 = isInit ? _GEN_7 : inputMemBound;
  assign _GEN_19 = isInit ? _GEN_14 : outputMemAddr;
  assign _GEN_20 = isInit ? _GEN_11 : outputLenAddr;
  assign _GEN_21 = isInit ? _GEN_12 : isInit;
  assign _GEN_22 = isInit ? _GEN_13 : initDone;
  assign _GEN_23 = io_inputMemBlockValid ? _GEN_16 : _GEN_1;
  assign _GEN_24 = io_inputMemBlockValid ? _GEN_17 : inputBitsRemaining;
  assign _GEN_25 = io_inputMemBlockValid ? _GEN_18 : inputMemBound;
  assign _GEN_26 = io_inputMemBlockValid ? _GEN_19 : outputMemAddr;
  assign _GEN_27 = io_inputMemBlockValid ? _GEN_20 : outputLenAddr;
  assign _GEN_28 = io_inputMemBlockValid ? _GEN_21 : isInit;
  assign _GEN_29 = io_inputMemBlockValid ? _GEN_22 : initDone;
  assign _T_139 = core_io_inputMemConsumed & _T_58;
  assign _GEN_30 = _T_139 ? 1'h1 : coreInputFinished;
  assign _GEN_31 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_146 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_148 = outputAddressAccepted == 1'h0;
  assign _T_150 = outputLengthCommitted == 1'h0;
  assign _T_151 = core_io_outputFinished & _T_150;
  assign _T_152 = core_io_outputMemBlockValid | _T_151;
  assign _T_153 = _T_148 & _T_152;
  assign _T_154 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _GEN_32 = _T_154 ? 1'h1 : outputAddressAccepted;
  assign _T_160 = outputBlockCounter == 5'h1f;
  assign _GEN_33 = io_outputMemBlockReady ? 5'h0 : outputBlockCounter;
  assign _T_163 = outputBlockCounter + 5'h1;
  assign _T_164 = _T_163[4:0];
  assign _GEN_34 = _T_160 ? _GEN_33 : _T_164;
  assign _GEN_35 = outputAddressAcceptedNext ? _GEN_34 : outputBlockCounter;
  assign _T_167 = outputBlockCounter == 5'h0;
  assign _T_168 = outputBits[15:0];
  assign _T_170 = outputBlockCounter == 5'h1;
  assign _T_171 = outputBits[31:16];
  assign _T_173 = _T_170 ? _T_171 : 16'h0;
  assign _T_174 = _T_167 ? _T_168 : _T_173;
  assign _T_175 = core_io_outputFinished ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_176 = outputAddressAcceptedNext & io_outputMemBlockReady;
  assign _T_180 = _T_176 & _T_160;
  assign _GEN_48 = {{22'd0}, core_io_outputBits};
  assign _T_184 = outputBits + _GEN_48;
  assign _T_185 = _T_184[31:0];
  assign _GEN_36 = core_io_outputFinished ? 1'h1 : outputLengthCommitted;
  assign _GEN_37 = core_io_outputFinished ? outputBits : _T_185;
  assign _GEN_38 = core_io_outputFinished ? _GEN_26 : _T_124;
  assign _GEN_39 = _T_180 ? 1'h0 : _GEN_32;
  assign _GEN_40 = _T_180 ? 1'h0 : _GEN_31;
  assign _GEN_41 = _T_180 ? _GEN_36 : outputLengthCommitted;
  assign _GEN_42 = _T_180 ? _GEN_37 : outputBits;
  assign _GEN_43 = _T_180 ? _GEN_38 : _GEN_26;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemBlockReady = _T_62;
  assign io_outputMemAddr = _T_146;
  assign io_outputMemAddrValid = _T_153;
  assign io_outputMemBlock = _T_175;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_inputAddrsIgnore = _T_55;
  assign io_inputBlocksFinished = _T_58;
  assign io_outputFinished = outputLengthCommitted;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_63;
  assign core_io_inputBits = _T_67[9:0];
  assign core_io_inputFinished = coreInputFinished;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_io_outputMemFlushed = _T_176;
  assign core_clock = clock;
  assign core_reset = reset;
  assign outputBitsBlock = _T_174;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputBitsRemaining = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  coreInputFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  outputBits = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputBlockCounter = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputLengthCommitted = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemAddr = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBound = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  outputMemAddr = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  outputLenAddr = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  initAddressAcked = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  outputAddressAccepted = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  outputAddressAcceptedNext = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_119) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_119) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 32'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_94) begin
            inputBitsRemaining <= _T_96;
          end else begin
            if (_T_77) begin
              inputBitsRemaining <= _T_79;
            end
          end
        end else begin
          if (_T_119) begin
            if (_T_65) begin
              inputBitsRemaining <= _T_132;
            end else begin
              inputBitsRemaining <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      coreInputFinished <= 1'h0;
    end else begin
      if (_T_139) begin
        coreInputFinished <= 1'h1;
      end
    end
    if (reset) begin
      outputBits <= 32'h0;
    end else begin
      if (_T_180) begin
        if (!(core_io_outputFinished)) begin
          outputBits <= _T_185;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_160) begin
          if (io_outputMemBlockReady) begin
            outputBlockCounter <= 5'h0;
          end
        end else begin
          outputBlockCounter <= _T_164;
        end
      end
    end
    if (reset) begin
      outputLengthCommitted <= 1'h0;
    end else begin
      if (_T_180) begin
        if (core_io_outputFinished) begin
          outputLengthCommitted <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= 32'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_73) begin
            inputMemAddr <= _T_75;
          end else begin
            if (_T_69) begin
              inputMemAddr <= _T_71;
            end else begin
              if (_T_48) begin
                inputMemAddr <= _T_51;
              end
            end
          end
        end else begin
          if (_T_48) begin
            inputMemAddr <= _T_51;
          end
        end
      end else begin
        if (_T_48) begin
          inputMemAddr <= _T_51;
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_94) begin
          inputMemBound <= _T_109;
        end else begin
          if (_T_77) begin
            inputMemBound <= _T_92;
          end
        end
      end
    end
    if (_T_180) begin
      if (core_io_outputFinished) begin
        if (io_inputMemBlockValid) begin
          if (isInit) begin
            if (_T_119) begin
              outputMemAddr <= _T_124;
            end else begin
              if (_T_115) begin
                outputMemAddr <= _T_117;
              end else begin
                if (_T_111) begin
                  outputMemAddr <= _T_113;
                end
              end
            end
          end
        end
      end else begin
        outputMemAddr <= _T_124;
      end
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_119) begin
            outputMemAddr <= _T_124;
          end else begin
            if (_T_115) begin
              outputMemAddr <= _T_117;
            end else begin
              if (_T_111) begin
                outputMemAddr <= _T_113;
              end
            end
          end
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_115) begin
          outputLenAddr <= _T_117;
        end else begin
          if (_T_111) begin
            outputLenAddr <= _T_113;
          end
        end
      end
    end
    if (reset) begin
      initAddressAcked <= 1'h0;
    end else begin
      if (io_inputMemAddrConsumed) begin
        initAddressAcked <= 1'h1;
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_180) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_154) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_180) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41 & _T_44) begin
          $fwrite(32'h80000002,"input address 0x%h accepted for core 1\n",io_inputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_154 & _T_44) begin
          $fwrite(32'h80000002,"output address 0x%h accepted for core 1\n",io_outputMemAddr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module StreamingWrapper(
  input          clock,
  input          reset,
  output [63:0]  io_inputMemAddrs_0,
  output [63:0]  io_inputMemAddrs_1,
  output         io_inputMemAddrValids_0,
  output         io_inputMemAddrValids_1,
  input          io_inputMemAddrReadys_0,
  input          io_inputMemAddrReadys_1,
  input  [511:0] io_inputMemBlocks_0,
  input  [511:0] io_inputMemBlocks_1,
  input          io_inputMemBlockValids_0,
  input          io_inputMemBlockValids_1,
  output         io_inputMemBlockReadys_0,
  output         io_inputMemBlockReadys_1,
  output [63:0]  io_outputMemAddrs_0,
  output [63:0]  io_outputMemAddrs_1,
  output         io_outputMemAddrValids_0,
  output         io_outputMemAddrValids_1,
  input          io_outputMemAddrReadys_0,
  input          io_outputMemAddrReadys_1,
  output [511:0] io_outputMemBlocks_0,
  output [511:0] io_outputMemBlocks_1,
  output         io_outputMemBlockValids_0,
  output         io_outputMemBlockValids_1,
  input          io_outputMemBlockReadys_0,
  input          io_outputMemBlockReadys_1,
  output         io_finished
);
  wire  StreamingCore_clock;
  wire  StreamingCore_reset;
  wire [31:0] StreamingCore_io_inputMemAddr;
  wire  StreamingCore_io_inputMemAddrConsumed;
  wire [15:0] StreamingCore_io_inputMemBlock;
  wire [4:0] StreamingCore_io_inputMemIdx;
  wire  StreamingCore_io_inputMemBlockValid;
  wire  StreamingCore_io_inputMemBlockReady;
  wire [31:0] StreamingCore_io_outputMemAddr;
  wire  StreamingCore_io_outputMemAddrValid;
  wire  StreamingCore_io_outputMemAddrReady;
  wire [15:0] StreamingCore_io_outputMemBlock;
  wire [4:0] StreamingCore_io_outputMemIdx;
  wire  StreamingCore_io_outputMemBlockValid;
  wire  StreamingCore_io_outputMemBlockReady;
  wire  StreamingCore_io_inputAddrsIgnore;
  wire  StreamingCore_io_inputBlocksFinished;
  wire  StreamingCore_io_outputFinished;
  wire  StreamingCore_1_clock;
  wire  StreamingCore_1_reset;
  wire [31:0] StreamingCore_1_io_inputMemAddr;
  wire  StreamingCore_1_io_inputMemAddrConsumed;
  wire [15:0] StreamingCore_1_io_inputMemBlock;
  wire [4:0] StreamingCore_1_io_inputMemIdx;
  wire  StreamingCore_1_io_inputMemBlockValid;
  wire  StreamingCore_1_io_inputMemBlockReady;
  wire [31:0] StreamingCore_1_io_outputMemAddr;
  wire  StreamingCore_1_io_outputMemAddrValid;
  wire  StreamingCore_1_io_outputMemAddrReady;
  wire [15:0] StreamingCore_1_io_outputMemBlock;
  wire [4:0] StreamingCore_1_io_outputMemIdx;
  wire  StreamingCore_1_io_outputMemBlockValid;
  wire  StreamingCore_1_io_outputMemBlockReady;
  wire  StreamingCore_1_io_inputAddrsIgnore;
  wire  StreamingCore_1_io_inputBlocksFinished;
  wire  StreamingCore_1_io_outputFinished;
  wire [31:0] cores_0_inputMemAddr;
  wire  cores_0_inputMemAddrConsumed;
  wire [15:0] cores_0_inputMemBlock;
  wire [4:0] cores_0_inputMemIdx;
  wire  cores_0_inputMemBlockValid;
  wire  cores_0_inputMemBlockReady;
  wire [31:0] cores_0_outputMemAddr;
  wire  cores_0_outputMemAddrValid;
  wire  cores_0_outputMemAddrReady;
  wire [15:0] cores_0_outputMemBlock;
  wire [4:0] cores_0_outputMemIdx;
  wire  cores_0_outputMemBlockValid;
  wire  cores_0_outputMemBlockReady;
  wire  cores_0_inputAddrsIgnore;
  wire  cores_0_inputBlocksFinished;
  wire  cores_0_outputFinished;
  wire [31:0] cores_1_inputMemAddr;
  wire  cores_1_inputMemAddrConsumed;
  wire [15:0] cores_1_inputMemBlock;
  wire [4:0] cores_1_inputMemIdx;
  wire  cores_1_inputMemBlockValid;
  wire  cores_1_inputMemBlockReady;
  wire [31:0] cores_1_outputMemAddr;
  wire  cores_1_outputMemAddrValid;
  wire  cores_1_outputMemAddrReady;
  wire [15:0] cores_1_outputMemBlock;
  wire [4:0] cores_1_outputMemIdx;
  wire  cores_1_outputMemBlockValid;
  wire  cores_1_outputMemBlockReady;
  wire  cores_1_inputAddrsIgnore;
  wire  cores_1_inputBlocksFinished;
  wire  cores_1_outputFinished;
  reg  _T_239;
  reg [31:0] _RAND_0;
  reg  _T_242;
  reg [31:0] _RAND_1;
  reg  _T_245;
  reg [31:0] _RAND_2;
  reg  _T_248;
  reg [31:0] _RAND_3;
  reg  _T_251;
  reg [31:0] _RAND_4;
  reg  _T_254;
  reg [31:0] _RAND_5;
  reg [31:0] _T_256;
  reg [31:0] _RAND_6;
  reg  _T_258;
  reg [31:0] _RAND_7;
  reg  _T_260;
  reg [31:0] _RAND_8;
  reg  _T_262;
  reg [31:0] _RAND_9;
  wire [31:0] _T_265_0;
  wire  _T_271_0;
  wire  _T_277_0;
  wire  _T_283_0;
  reg [31:0] _T_288;
  reg [31:0] _RAND_10;
  reg  _T_290;
  reg [31:0] _RAND_11;
  reg  _T_292;
  reg [31:0] _RAND_12;
  reg  _T_294;
  reg [31:0] _RAND_13;
  wire [31:0] _T_297_0;
  wire  _T_303_0;
  wire  _T_309_0;
  wire  _T_315_0;
  reg [31:0] _T_320;
  reg [31:0] _RAND_14;
  reg  _T_322;
  reg [31:0] _RAND_15;
  reg  _T_324;
  reg [31:0] _RAND_16;
  reg [15:0] _T_326;
  reg [31:0] _RAND_17;
  reg [4:0] _T_328;
  reg [31:0] _RAND_18;
  reg  _T_330;
  reg [31:0] _RAND_19;
  wire [31:0] _T_333_0;
  wire  _T_339_0;
  wire  _T_345_0;
  wire [15:0] _T_351_0;
  wire [4:0] _T_357_0;
  wire  _T_363_0;
  reg [31:0] _T_368;
  reg [31:0] _RAND_20;
  reg  _T_370;
  reg [31:0] _RAND_21;
  reg  _T_372;
  reg [31:0] _RAND_22;
  reg [15:0] _T_374;
  reg [31:0] _RAND_23;
  reg [4:0] _T_376;
  reg [31:0] _RAND_24;
  reg  _T_378;
  reg [31:0] _RAND_25;
  wire [31:0] _T_381_0;
  wire  _T_387_0;
  wire  _T_393_0;
  wire [15:0] _T_399_0;
  wire [4:0] _T_405_0;
  wire  _T_411_0;
  reg  _T_417;
  reg [31:0] _RAND_26;
  wire  _T_419;
  wire [1:0] _T_421;
  wire  _T_422;
  wire  _GEN_4;
  reg  _T_425;
  reg [31:0] _RAND_27;
  wire  _T_430;
  wire  _T_431;
  wire  _T_433;
  wire  _T_435;
  wire [1:0] _T_438;
  wire  _T_439;
  wire  _T_440;
  wire [1:0] _T_444;
  wire  _T_445;
  wire  _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _T_453;
  wire  _T_454;
  reg  _T_457;
  reg [31:0] _RAND_28;
  wire  _T_459;
  wire [1:0] _T_461;
  wire  _T_462;
  wire  _GEN_11;
  reg [15:0] _T_536_0_0;
  reg [31:0] _RAND_29;
  reg [15:0] _T_536_0_1;
  reg [31:0] _RAND_30;
  reg [15:0] _T_536_0_2;
  reg [31:0] _RAND_31;
  reg [15:0] _T_536_0_3;
  reg [31:0] _RAND_32;
  reg [15:0] _T_536_0_4;
  reg [31:0] _RAND_33;
  reg [15:0] _T_536_0_5;
  reg [31:0] _RAND_34;
  reg [15:0] _T_536_0_6;
  reg [31:0] _RAND_35;
  reg [15:0] _T_536_0_7;
  reg [31:0] _RAND_36;
  reg [15:0] _T_536_0_8;
  reg [31:0] _RAND_37;
  reg [15:0] _T_536_0_9;
  reg [31:0] _RAND_38;
  reg [15:0] _T_536_0_10;
  reg [31:0] _RAND_39;
  reg [15:0] _T_536_0_11;
  reg [31:0] _RAND_40;
  reg [15:0] _T_536_0_12;
  reg [31:0] _RAND_41;
  reg [15:0] _T_536_0_13;
  reg [31:0] _RAND_42;
  reg [15:0] _T_536_0_14;
  reg [31:0] _RAND_43;
  reg [15:0] _T_536_0_15;
  reg [31:0] _RAND_44;
  reg [15:0] _T_536_0_16;
  reg [31:0] _RAND_45;
  reg [15:0] _T_536_0_17;
  reg [31:0] _RAND_46;
  reg [15:0] _T_536_0_18;
  reg [31:0] _RAND_47;
  reg [15:0] _T_536_0_19;
  reg [31:0] _RAND_48;
  reg [15:0] _T_536_0_20;
  reg [31:0] _RAND_49;
  reg [15:0] _T_536_0_21;
  reg [31:0] _RAND_50;
  reg [15:0] _T_536_0_22;
  reg [31:0] _RAND_51;
  reg [15:0] _T_536_0_23;
  reg [31:0] _RAND_52;
  reg [15:0] _T_536_0_24;
  reg [31:0] _RAND_53;
  reg [15:0] _T_536_0_25;
  reg [31:0] _RAND_54;
  reg [15:0] _T_536_0_26;
  reg [31:0] _RAND_55;
  reg [15:0] _T_536_0_27;
  reg [31:0] _RAND_56;
  reg [15:0] _T_536_0_28;
  reg [31:0] _RAND_57;
  reg [15:0] _T_536_0_29;
  reg [31:0] _RAND_58;
  reg [15:0] _T_536_0_30;
  reg [31:0] _RAND_59;
  reg [15:0] _T_536_0_31;
  reg [31:0] _RAND_60;
  reg [4:0] _T_755_0;
  reg [31:0] _RAND_61;
  reg  _T_776_0;
  reg [31:0] _RAND_62;
  reg  _T_786;
  reg [31:0] _RAND_63;
  wire  _T_792;
  wire  _T_793;
  wire  _T_794;
  wire  _T_797;
  wire  _T_798;
  wire [15:0] _T_902;
  wire [15:0] _T_1006;
  wire [15:0] _T_1110;
  wire [15:0] _T_1214;
  wire [15:0] _T_1318;
  wire [15:0] _T_1422;
  wire [15:0] _T_1526;
  wire [15:0] _T_1630;
  wire [15:0] _T_1734;
  wire [15:0] _T_1838;
  wire [15:0] _T_1942;
  wire [15:0] _T_2046;
  wire [15:0] _T_2150;
  wire [15:0] _T_2254;
  wire [15:0] _T_2358;
  wire [15:0] _T_2462;
  wire [15:0] _T_2566;
  wire [15:0] _T_2670;
  wire [15:0] _T_2774;
  wire [15:0] _T_2878;
  wire [15:0] _T_2982;
  wire [15:0] _T_3086;
  wire [15:0] _T_3190;
  wire [15:0] _T_3294;
  wire [15:0] _T_3398;
  wire [15:0] _T_3502;
  wire [15:0] _T_3606;
  wire [15:0] _T_3710;
  wire [15:0] _T_3814;
  wire [15:0] _T_3918;
  wire [15:0] _T_4022;
  wire [15:0] _T_4126;
  wire  _T_4134;
  wire [1:0] _T_4136;
  wire  _T_4137;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_15;
  wire [15:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [15:0] _GEN_20;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_22;
  wire [15:0] _GEN_23;
  wire [15:0] _GEN_24;
  wire [15:0] _GEN_25;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  wire [15:0] _GEN_32;
  wire [15:0] _GEN_33;
  wire [15:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire [15:0] _GEN_36;
  wire [15:0] _GEN_37;
  wire [15:0] _GEN_38;
  wire [15:0] _GEN_39;
  wire [15:0] _GEN_40;
  wire [15:0] _GEN_41;
  wire [15:0] _GEN_42;
  wire [15:0] _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _T_4141;
  wire  _T_4142;
  wire  _T_4144;
  wire [1:0] _T_4147;
  wire  _T_4148;
  wire  _T_4149;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire [1:0] _T_4153;
  wire  _T_4156;
  wire  _T_4158;
  wire [5:0] _T_4162;
  wire [4:0] _T_4163;
  wire  _GEN_49;
  wire [4:0] _GEN_50;
  wire  _GEN_51;
  wire [4:0] _GEN_52;
  wire  _T_4173;
  wire  _T_4178;
  wire  _T_4183;
  wire  _T_4184;
  wire  _T_4186;
  wire [15:0] _GEN_0;
  wire [15:0] _GEN_53;
  wire [15:0] _GEN_54;
  wire [15:0] _GEN_55;
  wire [15:0] _GEN_56;
  wire [15:0] _GEN_57;
  wire [15:0] _GEN_58;
  wire [15:0] _GEN_59;
  wire [15:0] _GEN_60;
  wire [15:0] _GEN_61;
  wire [15:0] _GEN_62;
  wire [15:0] _GEN_63;
  wire [15:0] _GEN_64;
  wire [15:0] _GEN_65;
  wire [15:0] _GEN_66;
  wire [15:0] _GEN_67;
  wire [15:0] _GEN_68;
  wire [15:0] _GEN_69;
  wire [15:0] _GEN_70;
  wire [15:0] _GEN_71;
  wire [15:0] _GEN_72;
  wire [15:0] _GEN_73;
  wire [15:0] _GEN_74;
  wire [15:0] _GEN_75;
  wire [15:0] _GEN_76;
  wire [15:0] _GEN_77;
  wire [15:0] _GEN_78;
  wire [15:0] _GEN_79;
  wire [15:0] _GEN_80;
  wire [15:0] _GEN_81;
  wire [15:0] _GEN_82;
  wire [15:0] _GEN_83;
  wire  _T_4192;
  reg  _T_4195;
  reg [31:0] _RAND_64;
  wire  _T_4197;
  wire [1:0] _T_4199;
  wire  _T_4200;
  wire  _GEN_84;
  reg  _T_4203;
  reg [31:0] _RAND_65;
  wire  _T_4208;
  wire  _T_4209;
  wire  _T_4211;
  wire [1:0] _T_4216;
  wire  _T_4217;
  wire  _T_4218;
  wire [1:0] _T_4222;
  wire  _T_4223;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire  _GEN_90;
  wire  _T_4231;
  wire  _T_4232;
  reg  _T_4235;
  reg [31:0] _RAND_66;
  wire  _T_4237;
  wire [1:0] _T_4239;
  wire  _T_4240;
  wire  _GEN_91;
  reg [15:0] _T_4314_0_0;
  reg [31:0] _RAND_67;
  reg [15:0] _T_4314_0_1;
  reg [31:0] _RAND_68;
  reg [15:0] _T_4314_0_2;
  reg [31:0] _RAND_69;
  reg [15:0] _T_4314_0_3;
  reg [31:0] _RAND_70;
  reg [15:0] _T_4314_0_4;
  reg [31:0] _RAND_71;
  reg [15:0] _T_4314_0_5;
  reg [31:0] _RAND_72;
  reg [15:0] _T_4314_0_6;
  reg [31:0] _RAND_73;
  reg [15:0] _T_4314_0_7;
  reg [31:0] _RAND_74;
  reg [15:0] _T_4314_0_8;
  reg [31:0] _RAND_75;
  reg [15:0] _T_4314_0_9;
  reg [31:0] _RAND_76;
  reg [15:0] _T_4314_0_10;
  reg [31:0] _RAND_77;
  reg [15:0] _T_4314_0_11;
  reg [31:0] _RAND_78;
  reg [15:0] _T_4314_0_12;
  reg [31:0] _RAND_79;
  reg [15:0] _T_4314_0_13;
  reg [31:0] _RAND_80;
  reg [15:0] _T_4314_0_14;
  reg [31:0] _RAND_81;
  reg [15:0] _T_4314_0_15;
  reg [31:0] _RAND_82;
  reg [15:0] _T_4314_0_16;
  reg [31:0] _RAND_83;
  reg [15:0] _T_4314_0_17;
  reg [31:0] _RAND_84;
  reg [15:0] _T_4314_0_18;
  reg [31:0] _RAND_85;
  reg [15:0] _T_4314_0_19;
  reg [31:0] _RAND_86;
  reg [15:0] _T_4314_0_20;
  reg [31:0] _RAND_87;
  reg [15:0] _T_4314_0_21;
  reg [31:0] _RAND_88;
  reg [15:0] _T_4314_0_22;
  reg [31:0] _RAND_89;
  reg [15:0] _T_4314_0_23;
  reg [31:0] _RAND_90;
  reg [15:0] _T_4314_0_24;
  reg [31:0] _RAND_91;
  reg [15:0] _T_4314_0_25;
  reg [31:0] _RAND_92;
  reg [15:0] _T_4314_0_26;
  reg [31:0] _RAND_93;
  reg [15:0] _T_4314_0_27;
  reg [31:0] _RAND_94;
  reg [15:0] _T_4314_0_28;
  reg [31:0] _RAND_95;
  reg [15:0] _T_4314_0_29;
  reg [31:0] _RAND_96;
  reg [15:0] _T_4314_0_30;
  reg [31:0] _RAND_97;
  reg [15:0] _T_4314_0_31;
  reg [31:0] _RAND_98;
  reg [4:0] _T_4533_0;
  reg [31:0] _RAND_99;
  reg  _T_4554_0;
  reg [31:0] _RAND_100;
  reg  _T_4564;
  reg [31:0] _RAND_101;
  wire  _T_4570;
  wire  _T_4571;
  wire  _T_4572;
  wire  _T_4575;
  wire  _T_4576;
  wire [15:0] _T_4680;
  wire [15:0] _T_4784;
  wire [15:0] _T_4888;
  wire [15:0] _T_4992;
  wire [15:0] _T_5096;
  wire [15:0] _T_5200;
  wire [15:0] _T_5304;
  wire [15:0] _T_5408;
  wire [15:0] _T_5512;
  wire [15:0] _T_5616;
  wire [15:0] _T_5720;
  wire [15:0] _T_5824;
  wire [15:0] _T_5928;
  wire [15:0] _T_6032;
  wire [15:0] _T_6136;
  wire [15:0] _T_6240;
  wire [15:0] _T_6344;
  wire [15:0] _T_6448;
  wire [15:0] _T_6552;
  wire [15:0] _T_6656;
  wire [15:0] _T_6760;
  wire [15:0] _T_6864;
  wire [15:0] _T_6968;
  wire [15:0] _T_7072;
  wire [15:0] _T_7176;
  wire [15:0] _T_7280;
  wire [15:0] _T_7384;
  wire [15:0] _T_7488;
  wire [15:0] _T_7592;
  wire [15:0] _T_7696;
  wire [15:0] _T_7800;
  wire [15:0] _T_7904;
  wire  _T_7912;
  wire [1:0] _T_7914;
  wire  _T_7915;
  wire [15:0] _GEN_92;
  wire [15:0] _GEN_93;
  wire [15:0] _GEN_94;
  wire [15:0] _GEN_95;
  wire [15:0] _GEN_96;
  wire [15:0] _GEN_97;
  wire [15:0] _GEN_98;
  wire [15:0] _GEN_99;
  wire [15:0] _GEN_100;
  wire [15:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire [15:0] _GEN_103;
  wire [15:0] _GEN_104;
  wire [15:0] _GEN_105;
  wire [15:0] _GEN_106;
  wire [15:0] _GEN_107;
  wire [15:0] _GEN_108;
  wire [15:0] _GEN_109;
  wire [15:0] _GEN_110;
  wire [15:0] _GEN_111;
  wire [15:0] _GEN_112;
  wire [15:0] _GEN_113;
  wire [15:0] _GEN_114;
  wire [15:0] _GEN_115;
  wire [15:0] _GEN_116;
  wire [15:0] _GEN_117;
  wire [15:0] _GEN_118;
  wire [15:0] _GEN_119;
  wire [15:0] _GEN_120;
  wire [15:0] _GEN_121;
  wire [15:0] _GEN_122;
  wire [15:0] _GEN_123;
  wire  _GEN_124;
  wire  _GEN_125;
  wire  _T_7919;
  wire  _T_7920;
  wire [1:0] _T_7925;
  wire  _T_7926;
  wire  _T_7927;
  wire  _GEN_126;
  wire  _GEN_127;
  wire  _GEN_128;
  wire [1:0] _T_7931;
  wire  _T_7936;
  wire [5:0] _T_7940;
  wire [4:0] _T_7941;
  wire  _GEN_129;
  wire [4:0] _GEN_130;
  wire  _GEN_131;
  wire [4:0] _GEN_132;
  wire  _T_7951;
  wire  _T_7956;
  wire  _T_7961;
  wire  _T_7962;
  wire  _T_7964;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_133;
  wire [15:0] _GEN_134;
  wire [15:0] _GEN_135;
  wire [15:0] _GEN_136;
  wire [15:0] _GEN_137;
  wire [15:0] _GEN_138;
  wire [15:0] _GEN_139;
  wire [15:0] _GEN_140;
  wire [15:0] _GEN_141;
  wire [15:0] _GEN_142;
  wire [15:0] _GEN_143;
  wire [15:0] _GEN_144;
  wire [15:0] _GEN_145;
  wire [15:0] _GEN_146;
  wire [15:0] _GEN_147;
  wire [15:0] _GEN_148;
  wire [15:0] _GEN_149;
  wire [15:0] _GEN_150;
  wire [15:0] _GEN_151;
  wire [15:0] _GEN_152;
  wire [15:0] _GEN_153;
  wire [15:0] _GEN_154;
  wire [15:0] _GEN_155;
  wire [15:0] _GEN_156;
  wire [15:0] _GEN_157;
  wire [15:0] _GEN_158;
  wire [15:0] _GEN_159;
  wire [15:0] _GEN_160;
  wire [15:0] _GEN_161;
  wire [15:0] _GEN_162;
  wire [15:0] _GEN_163;
  wire  _T_7970;
  reg  _T_7973;
  reg [31:0] _RAND_102;
  wire  _T_7975;
  wire [1:0] _T_7977;
  wire  _T_7978;
  wire  _GEN_164;
  reg  _T_7992_0;
  reg [31:0] _RAND_103;
  reg [31:0] _T_8003_0;
  reg [31:0] _RAND_104;
  reg [15:0] _T_8080_0_0;
  reg [31:0] _RAND_105;
  reg [15:0] _T_8080_0_1;
  reg [31:0] _RAND_106;
  reg [15:0] _T_8080_0_2;
  reg [31:0] _RAND_107;
  reg [15:0] _T_8080_0_3;
  reg [31:0] _RAND_108;
  reg [15:0] _T_8080_0_4;
  reg [31:0] _RAND_109;
  reg [15:0] _T_8080_0_5;
  reg [31:0] _RAND_110;
  reg [15:0] _T_8080_0_6;
  reg [31:0] _RAND_111;
  reg [15:0] _T_8080_0_7;
  reg [31:0] _RAND_112;
  reg [15:0] _T_8080_0_8;
  reg [31:0] _RAND_113;
  reg [15:0] _T_8080_0_9;
  reg [31:0] _RAND_114;
  reg [15:0] _T_8080_0_10;
  reg [31:0] _RAND_115;
  reg [15:0] _T_8080_0_11;
  reg [31:0] _RAND_116;
  reg [15:0] _T_8080_0_12;
  reg [31:0] _RAND_117;
  reg [15:0] _T_8080_0_13;
  reg [31:0] _RAND_118;
  reg [15:0] _T_8080_0_14;
  reg [31:0] _RAND_119;
  reg [15:0] _T_8080_0_15;
  reg [31:0] _RAND_120;
  reg [15:0] _T_8080_0_16;
  reg [31:0] _RAND_121;
  reg [15:0] _T_8080_0_17;
  reg [31:0] _RAND_122;
  reg [15:0] _T_8080_0_18;
  reg [31:0] _RAND_123;
  reg [15:0] _T_8080_0_19;
  reg [31:0] _RAND_124;
  reg [15:0] _T_8080_0_20;
  reg [31:0] _RAND_125;
  reg [15:0] _T_8080_0_21;
  reg [31:0] _RAND_126;
  reg [15:0] _T_8080_0_22;
  reg [31:0] _RAND_127;
  reg [15:0] _T_8080_0_23;
  reg [31:0] _RAND_128;
  reg [15:0] _T_8080_0_24;
  reg [31:0] _RAND_129;
  reg [15:0] _T_8080_0_25;
  reg [31:0] _RAND_130;
  reg [15:0] _T_8080_0_26;
  reg [31:0] _RAND_131;
  reg [15:0] _T_8080_0_27;
  reg [31:0] _RAND_132;
  reg [15:0] _T_8080_0_28;
  reg [31:0] _RAND_133;
  reg [15:0] _T_8080_0_29;
  reg [31:0] _RAND_134;
  reg [15:0] _T_8080_0_30;
  reg [31:0] _RAND_135;
  reg [15:0] _T_8080_0_31;
  reg [31:0] _RAND_136;
  reg  _T_8299_0;
  reg [31:0] _RAND_137;
  reg  _T_8309;
  reg [31:0] _RAND_138;
  reg  _T_8312;
  reg [31:0] _RAND_139;
  reg  _T_8315;
  reg [31:0] _RAND_140;
  wire  _T_8319;
  wire  _T_8320;
  wire  _GEN_165;
  wire  _T_8324;
  wire  _T_8326;
  wire  _T_8327;
  wire  _GEN_166;
  wire [15:0] _GEN_2;
  wire [15:0] _GEN_167;
  wire [15:0] _GEN_168;
  wire [15:0] _GEN_169;
  wire [15:0] _GEN_170;
  wire [15:0] _GEN_171;
  wire [15:0] _GEN_172;
  wire [15:0] _GEN_173;
  wire [15:0] _GEN_174;
  wire [15:0] _GEN_175;
  wire [15:0] _GEN_176;
  wire [15:0] _GEN_177;
  wire [15:0] _GEN_178;
  wire [15:0] _GEN_179;
  wire [15:0] _GEN_180;
  wire [15:0] _GEN_181;
  wire [15:0] _GEN_182;
  wire [15:0] _GEN_183;
  wire [15:0] _GEN_184;
  wire [15:0] _GEN_185;
  wire [15:0] _GEN_186;
  wire [15:0] _GEN_187;
  wire [15:0] _GEN_188;
  wire [15:0] _GEN_189;
  wire [15:0] _GEN_190;
  wire [15:0] _GEN_191;
  wire [15:0] _GEN_192;
  wire [15:0] _GEN_193;
  wire [15:0] _GEN_194;
  wire [15:0] _GEN_195;
  wire [15:0] _GEN_196;
  wire [15:0] _GEN_197;
  wire [15:0] _GEN_198;
  wire [15:0] _GEN_199;
  wire [15:0] _GEN_200;
  wire [15:0] _GEN_201;
  wire [15:0] _GEN_202;
  wire [15:0] _GEN_203;
  wire [15:0] _GEN_204;
  wire [15:0] _GEN_205;
  wire [15:0] _GEN_206;
  wire [15:0] _GEN_207;
  wire [15:0] _GEN_208;
  wire [15:0] _GEN_209;
  wire [15:0] _GEN_210;
  wire [15:0] _GEN_211;
  wire [15:0] _GEN_212;
  wire [15:0] _GEN_213;
  wire [15:0] _GEN_214;
  wire [15:0] _GEN_215;
  wire [15:0] _GEN_216;
  wire [15:0] _GEN_217;
  wire [15:0] _GEN_218;
  wire [15:0] _GEN_219;
  wire [15:0] _GEN_220;
  wire [15:0] _GEN_221;
  wire [15:0] _GEN_222;
  wire [15:0] _GEN_223;
  wire [15:0] _GEN_224;
  wire [15:0] _GEN_225;
  wire [15:0] _GEN_226;
  wire [15:0] _GEN_227;
  wire [15:0] _GEN_228;
  wire [15:0] _GEN_229;
  wire [15:0] _GEN_230;
  wire  _T_8333;
  wire  _T_8335;
  wire  _T_8336;
  wire  _T_8342;
  wire  _GEN_231;
  wire [31:0] _GEN_232;
  wire  _T_8351;
  wire  _T_8352;
  wire [31:0] _T_8456;
  wire [31:0] _T_8457;
  wire [63:0] _T_8458;
  wire [31:0] _T_8459;
  wire [31:0] _T_8460;
  wire [63:0] _T_8461;
  wire [127:0] _T_8462;
  wire [31:0] _T_8463;
  wire [31:0] _T_8464;
  wire [63:0] _T_8465;
  wire [31:0] _T_8466;
  wire [31:0] _T_8467;
  wire [63:0] _T_8468;
  wire [127:0] _T_8469;
  wire [255:0] _T_8470;
  wire [31:0] _T_8471;
  wire [31:0] _T_8472;
  wire [63:0] _T_8473;
  wire [31:0] _T_8474;
  wire [31:0] _T_8475;
  wire [63:0] _T_8476;
  wire [127:0] _T_8477;
  wire [31:0] _T_8478;
  wire [31:0] _T_8479;
  wire [63:0] _T_8480;
  wire [31:0] _T_8481;
  wire [31:0] _T_8482;
  wire [63:0] _T_8483;
  wire [127:0] _T_8484;
  wire [255:0] _T_8485;
  wire [511:0] _T_8486;
  wire  _T_8491;
  wire  _T_8493;
  wire  _T_8498;
  wire  _T_8501;
  wire  _T_8502;
  wire  _T_8509;
  wire  _T_8510;
  wire  _T_8511;
  wire  _GEN_233;
  wire  _T_8513;
  wire  _T_8514;
  wire  _T_8521;
  wire  _T_8522;
  wire  _T_8525;
  wire  _T_8527;
  wire [1:0] _T_8530;
  wire  _T_8531;
  wire  _T_8532;
  wire [1:0] _T_8539;
  wire  _T_8540;
  wire  _GEN_234;
  wire  _GEN_235;
  wire  _GEN_236;
  wire  _GEN_237;
  wire  _GEN_238;
  wire  _GEN_239;
  wire  _GEN_240;
  wire  _GEN_241;
  wire  _GEN_242;
  wire  _GEN_243;
  wire  _GEN_244;
  wire  _GEN_245;
  wire  _GEN_246;
  wire  _T_8556;
  wire  _T_8561;
  wire  _T_8562;
  wire  _T_8564;
  wire  _T_8565;
  wire [1:0] _T_8566;
  reg  _T_8572;
  reg [31:0] _RAND_141;
  wire  _T_8574;
  wire [1:0] _T_8576;
  wire  _T_8577;
  wire  _GEN_247;
  reg  _T_8591_0;
  reg [31:0] _RAND_142;
  reg [31:0] _T_8602_0;
  reg [31:0] _RAND_143;
  reg [15:0] _T_8679_0_0;
  reg [31:0] _RAND_144;
  reg [15:0] _T_8679_0_1;
  reg [31:0] _RAND_145;
  reg [15:0] _T_8679_0_2;
  reg [31:0] _RAND_146;
  reg [15:0] _T_8679_0_3;
  reg [31:0] _RAND_147;
  reg [15:0] _T_8679_0_4;
  reg [31:0] _RAND_148;
  reg [15:0] _T_8679_0_5;
  reg [31:0] _RAND_149;
  reg [15:0] _T_8679_0_6;
  reg [31:0] _RAND_150;
  reg [15:0] _T_8679_0_7;
  reg [31:0] _RAND_151;
  reg [15:0] _T_8679_0_8;
  reg [31:0] _RAND_152;
  reg [15:0] _T_8679_0_9;
  reg [31:0] _RAND_153;
  reg [15:0] _T_8679_0_10;
  reg [31:0] _RAND_154;
  reg [15:0] _T_8679_0_11;
  reg [31:0] _RAND_155;
  reg [15:0] _T_8679_0_12;
  reg [31:0] _RAND_156;
  reg [15:0] _T_8679_0_13;
  reg [31:0] _RAND_157;
  reg [15:0] _T_8679_0_14;
  reg [31:0] _RAND_158;
  reg [15:0] _T_8679_0_15;
  reg [31:0] _RAND_159;
  reg [15:0] _T_8679_0_16;
  reg [31:0] _RAND_160;
  reg [15:0] _T_8679_0_17;
  reg [31:0] _RAND_161;
  reg [15:0] _T_8679_0_18;
  reg [31:0] _RAND_162;
  reg [15:0] _T_8679_0_19;
  reg [31:0] _RAND_163;
  reg [15:0] _T_8679_0_20;
  reg [31:0] _RAND_164;
  reg [15:0] _T_8679_0_21;
  reg [31:0] _RAND_165;
  reg [15:0] _T_8679_0_22;
  reg [31:0] _RAND_166;
  reg [15:0] _T_8679_0_23;
  reg [31:0] _RAND_167;
  reg [15:0] _T_8679_0_24;
  reg [31:0] _RAND_168;
  reg [15:0] _T_8679_0_25;
  reg [31:0] _RAND_169;
  reg [15:0] _T_8679_0_26;
  reg [31:0] _RAND_170;
  reg [15:0] _T_8679_0_27;
  reg [31:0] _RAND_171;
  reg [15:0] _T_8679_0_28;
  reg [31:0] _RAND_172;
  reg [15:0] _T_8679_0_29;
  reg [31:0] _RAND_173;
  reg [15:0] _T_8679_0_30;
  reg [31:0] _RAND_174;
  reg [15:0] _T_8679_0_31;
  reg [31:0] _RAND_175;
  reg  _T_8898_0;
  reg [31:0] _RAND_176;
  reg  _T_8908;
  reg [31:0] _RAND_177;
  reg  _T_8911;
  reg [31:0] _RAND_178;
  reg  _T_8914;
  reg [31:0] _RAND_179;
  wire  _T_8918;
  wire  _T_8919;
  wire  _GEN_248;
  wire  _T_8923;
  wire  _T_8925;
  wire  _T_8926;
  wire  _GEN_249;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_250;
  wire [15:0] _GEN_251;
  wire [15:0] _GEN_252;
  wire [15:0] _GEN_253;
  wire [15:0] _GEN_254;
  wire [15:0] _GEN_255;
  wire [15:0] _GEN_256;
  wire [15:0] _GEN_257;
  wire [15:0] _GEN_258;
  wire [15:0] _GEN_259;
  wire [15:0] _GEN_260;
  wire [15:0] _GEN_261;
  wire [15:0] _GEN_262;
  wire [15:0] _GEN_263;
  wire [15:0] _GEN_264;
  wire [15:0] _GEN_265;
  wire [15:0] _GEN_266;
  wire [15:0] _GEN_267;
  wire [15:0] _GEN_268;
  wire [15:0] _GEN_269;
  wire [15:0] _GEN_270;
  wire [15:0] _GEN_271;
  wire [15:0] _GEN_272;
  wire [15:0] _GEN_273;
  wire [15:0] _GEN_274;
  wire [15:0] _GEN_275;
  wire [15:0] _GEN_276;
  wire [15:0] _GEN_277;
  wire [15:0] _GEN_278;
  wire [15:0] _GEN_279;
  wire [15:0] _GEN_280;
  wire [15:0] _GEN_281;
  wire [15:0] _GEN_282;
  wire [15:0] _GEN_283;
  wire [15:0] _GEN_284;
  wire [15:0] _GEN_285;
  wire [15:0] _GEN_286;
  wire [15:0] _GEN_287;
  wire [15:0] _GEN_288;
  wire [15:0] _GEN_289;
  wire [15:0] _GEN_290;
  wire [15:0] _GEN_291;
  wire [15:0] _GEN_292;
  wire [15:0] _GEN_293;
  wire [15:0] _GEN_294;
  wire [15:0] _GEN_295;
  wire [15:0] _GEN_296;
  wire [15:0] _GEN_297;
  wire [15:0] _GEN_298;
  wire [15:0] _GEN_299;
  wire [15:0] _GEN_300;
  wire [15:0] _GEN_301;
  wire [15:0] _GEN_302;
  wire [15:0] _GEN_303;
  wire [15:0] _GEN_304;
  wire [15:0] _GEN_305;
  wire [15:0] _GEN_306;
  wire [15:0] _GEN_307;
  wire [15:0] _GEN_308;
  wire [15:0] _GEN_309;
  wire [15:0] _GEN_310;
  wire [15:0] _GEN_311;
  wire [15:0] _GEN_312;
  wire [15:0] _GEN_313;
  wire  _T_8932;
  wire  _T_8934;
  wire  _T_8935;
  wire  _T_8941;
  wire  _GEN_314;
  wire [31:0] _GEN_315;
  wire  _T_8950;
  wire  _T_8951;
  wire [31:0] _T_9055;
  wire [31:0] _T_9056;
  wire [63:0] _T_9057;
  wire [31:0] _T_9058;
  wire [31:0] _T_9059;
  wire [63:0] _T_9060;
  wire [127:0] _T_9061;
  wire [31:0] _T_9062;
  wire [31:0] _T_9063;
  wire [63:0] _T_9064;
  wire [31:0] _T_9065;
  wire [31:0] _T_9066;
  wire [63:0] _T_9067;
  wire [127:0] _T_9068;
  wire [255:0] _T_9069;
  wire [31:0] _T_9070;
  wire [31:0] _T_9071;
  wire [63:0] _T_9072;
  wire [31:0] _T_9073;
  wire [31:0] _T_9074;
  wire [63:0] _T_9075;
  wire [127:0] _T_9076;
  wire [31:0] _T_9077;
  wire [31:0] _T_9078;
  wire [63:0] _T_9079;
  wire [31:0] _T_9080;
  wire [31:0] _T_9081;
  wire [63:0] _T_9082;
  wire [127:0] _T_9083;
  wire [255:0] _T_9084;
  wire [511:0] _T_9085;
  wire  _T_9090;
  wire  _T_9092;
  wire  _T_9097;
  wire  _T_9100;
  wire  _T_9101;
  wire  _T_9108;
  wire  _T_9109;
  wire  _T_9110;
  wire  _GEN_316;
  wire  _T_9112;
  wire  _T_9113;
  wire  _T_9120;
  wire  _T_9121;
  wire  _T_9124;
  wire [1:0] _T_9129;
  wire  _T_9130;
  wire  _T_9131;
  wire [1:0] _T_9138;
  wire  _T_9139;
  wire  _GEN_317;
  wire  _GEN_318;
  wire  _GEN_319;
  wire  _GEN_320;
  wire  _GEN_321;
  wire  _GEN_322;
  wire  _GEN_323;
  wire  _GEN_324;
  wire  _GEN_325;
  wire  _GEN_326;
  wire  _GEN_327;
  wire  _GEN_328;
  wire  _GEN_329;
  wire  _T_9155;
  wire  _T_9160;
  wire  _T_9161;
  wire  _T_9163;
  wire  _T_9164;
  wire [1:0] _T_9165;
  wire  cumFinished;
  StreamingCore StreamingCore (
    .clock(StreamingCore_clock),
    .reset(StreamingCore_reset),
    .io_inputMemAddr(StreamingCore_io_inputMemAddr),
    .io_inputMemAddrConsumed(StreamingCore_io_inputMemAddrConsumed),
    .io_inputMemBlock(StreamingCore_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_io_outputMemBlockReady),
    .io_inputAddrsIgnore(StreamingCore_io_inputAddrsIgnore),
    .io_inputBlocksFinished(StreamingCore_io_inputBlocksFinished),
    .io_outputFinished(StreamingCore_io_outputFinished)
  );
  StreamingCore_1 StreamingCore_1 (
    .clock(StreamingCore_1_clock),
    .reset(StreamingCore_1_reset),
    .io_inputMemAddr(StreamingCore_1_io_inputMemAddr),
    .io_inputMemAddrConsumed(StreamingCore_1_io_inputMemAddrConsumed),
    .io_inputMemBlock(StreamingCore_1_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_1_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_1_io_inputMemBlockValid),
    .io_inputMemBlockReady(StreamingCore_1_io_inputMemBlockReady),
    .io_outputMemAddr(StreamingCore_1_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_1_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_1_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_1_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_1_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_1_io_outputMemBlockValid),
    .io_outputMemBlockReady(StreamingCore_1_io_outputMemBlockReady),
    .io_inputAddrsIgnore(StreamingCore_1_io_inputAddrsIgnore),
    .io_inputBlocksFinished(StreamingCore_1_io_inputBlocksFinished),
    .io_outputFinished(StreamingCore_1_io_outputFinished)
  );
  assign _T_419 = _T_417 != 1'h1;
  assign _T_421 = _T_417 + 1'h1;
  assign _T_422 = _T_421[0:0];
  assign _GEN_4 = _T_419 ? _T_422 : _T_417;
  assign _T_430 = io_inputMemAddrReadys_0 | _T_277_0;
  assign _T_431 = _T_417 & _T_430;
  assign _T_433 = _T_425 == 1'h0;
  assign _T_435 = _T_239 == 1'h0;
  assign _T_438 = _T_239 + 1'h1;
  assign _T_439 = _T_438[0:0];
  assign _T_440 = _T_435 ? 1'h0 : _T_439;
  assign _T_444 = _T_425 + 1'h1;
  assign _T_445 = _T_444[0:0];
  assign _GEN_5 = _T_433 ? _T_440 : _T_239;
  assign _GEN_6 = _T_433 ? 1'h0 : _GEN_4;
  assign _GEN_7 = _T_433 ? 1'h0 : _T_445;
  assign _GEN_8 = _T_431 ? _GEN_5 : _T_239;
  assign _GEN_9 = _T_431 ? _GEN_6 : _GEN_4;
  assign _GEN_10 = _T_431 ? _GEN_7 : _T_425;
  assign _T_453 = _T_277_0 == 1'h0;
  assign _T_454 = _T_417 & _T_453;
  assign _T_459 = _T_457 != 1'h1;
  assign _T_461 = _T_457 + 1'h1;
  assign _T_462 = _T_461[0:0];
  assign _GEN_11 = _T_459 ? _T_462 : _T_457;
  assign _T_792 = _T_786 == 1'h0;
  assign _T_793 = _T_457 & _T_792;
  assign _T_794 = io_inputMemBlockReadys_0 & io_inputMemBlockValids_0;
  assign _T_797 = _T_794 | _T_283_0;
  assign _T_798 = _T_793 & _T_797;
  assign _T_902 = io_inputMemBlocks_0[15:0];
  assign _T_1006 = io_inputMemBlocks_0[31:16];
  assign _T_1110 = io_inputMemBlocks_0[47:32];
  assign _T_1214 = io_inputMemBlocks_0[63:48];
  assign _T_1318 = io_inputMemBlocks_0[79:64];
  assign _T_1422 = io_inputMemBlocks_0[95:80];
  assign _T_1526 = io_inputMemBlocks_0[111:96];
  assign _T_1630 = io_inputMemBlocks_0[127:112];
  assign _T_1734 = io_inputMemBlocks_0[143:128];
  assign _T_1838 = io_inputMemBlocks_0[159:144];
  assign _T_1942 = io_inputMemBlocks_0[175:160];
  assign _T_2046 = io_inputMemBlocks_0[191:176];
  assign _T_2150 = io_inputMemBlocks_0[207:192];
  assign _T_2254 = io_inputMemBlocks_0[223:208];
  assign _T_2358 = io_inputMemBlocks_0[239:224];
  assign _T_2462 = io_inputMemBlocks_0[255:240];
  assign _T_2566 = io_inputMemBlocks_0[271:256];
  assign _T_2670 = io_inputMemBlocks_0[287:272];
  assign _T_2774 = io_inputMemBlocks_0[303:288];
  assign _T_2878 = io_inputMemBlocks_0[319:304];
  assign _T_2982 = io_inputMemBlocks_0[335:320];
  assign _T_3086 = io_inputMemBlocks_0[351:336];
  assign _T_3190 = io_inputMemBlocks_0[367:352];
  assign _T_3294 = io_inputMemBlocks_0[383:368];
  assign _T_3398 = io_inputMemBlocks_0[399:384];
  assign _T_3502 = io_inputMemBlocks_0[415:400];
  assign _T_3606 = io_inputMemBlocks_0[431:416];
  assign _T_3710 = io_inputMemBlocks_0[447:432];
  assign _T_3814 = io_inputMemBlocks_0[463:448];
  assign _T_3918 = io_inputMemBlocks_0[479:464];
  assign _T_4022 = io_inputMemBlocks_0[495:480];
  assign _T_4126 = io_inputMemBlocks_0[511:496];
  assign _T_4134 = _T_283_0 == 1'h0;
  assign _T_4136 = _T_786 + 1'h1;
  assign _T_4137 = _T_4136[0:0];
  assign _GEN_12 = _T_798 ? _T_902 : _T_536_0_0;
  assign _GEN_13 = _T_798 ? _T_1006 : _T_536_0_1;
  assign _GEN_14 = _T_798 ? _T_1110 : _T_536_0_2;
  assign _GEN_15 = _T_798 ? _T_1214 : _T_536_0_3;
  assign _GEN_16 = _T_798 ? _T_1318 : _T_536_0_4;
  assign _GEN_17 = _T_798 ? _T_1422 : _T_536_0_5;
  assign _GEN_18 = _T_798 ? _T_1526 : _T_536_0_6;
  assign _GEN_19 = _T_798 ? _T_1630 : _T_536_0_7;
  assign _GEN_20 = _T_798 ? _T_1734 : _T_536_0_8;
  assign _GEN_21 = _T_798 ? _T_1838 : _T_536_0_9;
  assign _GEN_22 = _T_798 ? _T_1942 : _T_536_0_10;
  assign _GEN_23 = _T_798 ? _T_2046 : _T_536_0_11;
  assign _GEN_24 = _T_798 ? _T_2150 : _T_536_0_12;
  assign _GEN_25 = _T_798 ? _T_2254 : _T_536_0_13;
  assign _GEN_26 = _T_798 ? _T_2358 : _T_536_0_14;
  assign _GEN_27 = _T_798 ? _T_2462 : _T_536_0_15;
  assign _GEN_28 = _T_798 ? _T_2566 : _T_536_0_16;
  assign _GEN_29 = _T_798 ? _T_2670 : _T_536_0_17;
  assign _GEN_30 = _T_798 ? _T_2774 : _T_536_0_18;
  assign _GEN_31 = _T_798 ? _T_2878 : _T_536_0_19;
  assign _GEN_32 = _T_798 ? _T_2982 : _T_536_0_20;
  assign _GEN_33 = _T_798 ? _T_3086 : _T_536_0_21;
  assign _GEN_34 = _T_798 ? _T_3190 : _T_536_0_22;
  assign _GEN_35 = _T_798 ? _T_3294 : _T_536_0_23;
  assign _GEN_36 = _T_798 ? _T_3398 : _T_536_0_24;
  assign _GEN_37 = _T_798 ? _T_3502 : _T_536_0_25;
  assign _GEN_38 = _T_798 ? _T_3606 : _T_536_0_26;
  assign _GEN_39 = _T_798 ? _T_3710 : _T_536_0_27;
  assign _GEN_40 = _T_798 ? _T_3814 : _T_536_0_28;
  assign _GEN_41 = _T_798 ? _T_3918 : _T_536_0_29;
  assign _GEN_42 = _T_798 ? _T_4022 : _T_536_0_30;
  assign _GEN_43 = _T_798 ? _T_4126 : _T_536_0_31;
  assign _GEN_44 = _T_798 ? _T_4134 : _T_776_0;
  assign _GEN_45 = _T_798 ? _T_4137 : _T_786;
  assign _T_4141 = _T_776_0 == 1'h0;
  assign _T_4142 = _T_786 & _T_4141;
  assign _T_4144 = _T_242 == 1'h0;
  assign _T_4147 = _T_242 + 1'h1;
  assign _T_4148 = _T_4147[0:0];
  assign _T_4149 = _T_4144 ? 1'h0 : _T_4148;
  assign _GEN_46 = _T_4142 ? _T_4149 : _T_242;
  assign _GEN_47 = _T_4142 ? 1'h0 : _GEN_11;
  assign _GEN_48 = _T_4142 ? 1'h0 : _GEN_45;
  assign _T_4153 = {_T_242,_T_786};
  assign _T_4156 = reset == 1'h0;
  assign _T_4158 = _T_755_0 == 5'h1f;
  assign _T_4162 = _T_755_0 + 5'h1;
  assign _T_4163 = _T_4162[4:0];
  assign _GEN_49 = _T_4158 ? 1'h0 : _GEN_44;
  assign _GEN_50 = _T_4158 ? 5'h0 : _T_4163;
  assign _GEN_51 = _T_776_0 ? _GEN_49 : _GEN_44;
  assign _GEN_52 = _T_776_0 ? _GEN_50 : _T_755_0;
  assign _T_4173 = _T_793 & _T_271_0;
  assign _T_4178 = _T_4173 & _T_4134;
  assign _T_4183 = _T_433 & io_inputMemAddrReadys_0;
  assign _T_4184 = _T_4183 & io_inputMemAddrValids_0;
  assign _T_4186 = _T_435 ? _T_4184 : 1'h0;
  assign _GEN_53 = 5'h1 == _T_755_0 ? _T_536_0_1 : _T_536_0_0;
  assign _GEN_54 = 5'h2 == _T_755_0 ? _T_536_0_2 : _GEN_53;
  assign _GEN_55 = 5'h3 == _T_755_0 ? _T_536_0_3 : _GEN_54;
  assign _GEN_56 = 5'h4 == _T_755_0 ? _T_536_0_4 : _GEN_55;
  assign _GEN_57 = 5'h5 == _T_755_0 ? _T_536_0_5 : _GEN_56;
  assign _GEN_58 = 5'h6 == _T_755_0 ? _T_536_0_6 : _GEN_57;
  assign _GEN_59 = 5'h7 == _T_755_0 ? _T_536_0_7 : _GEN_58;
  assign _GEN_60 = 5'h8 == _T_755_0 ? _T_536_0_8 : _GEN_59;
  assign _GEN_61 = 5'h9 == _T_755_0 ? _T_536_0_9 : _GEN_60;
  assign _GEN_62 = 5'ha == _T_755_0 ? _T_536_0_10 : _GEN_61;
  assign _GEN_63 = 5'hb == _T_755_0 ? _T_536_0_11 : _GEN_62;
  assign _GEN_64 = 5'hc == _T_755_0 ? _T_536_0_12 : _GEN_63;
  assign _GEN_65 = 5'hd == _T_755_0 ? _T_536_0_13 : _GEN_64;
  assign _GEN_66 = 5'he == _T_755_0 ? _T_536_0_14 : _GEN_65;
  assign _GEN_67 = 5'hf == _T_755_0 ? _T_536_0_15 : _GEN_66;
  assign _GEN_68 = 5'h10 == _T_755_0 ? _T_536_0_16 : _GEN_67;
  assign _GEN_69 = 5'h11 == _T_755_0 ? _T_536_0_17 : _GEN_68;
  assign _GEN_70 = 5'h12 == _T_755_0 ? _T_536_0_18 : _GEN_69;
  assign _GEN_71 = 5'h13 == _T_755_0 ? _T_536_0_19 : _GEN_70;
  assign _GEN_72 = 5'h14 == _T_755_0 ? _T_536_0_20 : _GEN_71;
  assign _GEN_73 = 5'h15 == _T_755_0 ? _T_536_0_21 : _GEN_72;
  assign _GEN_74 = 5'h16 == _T_755_0 ? _T_536_0_22 : _GEN_73;
  assign _GEN_75 = 5'h17 == _T_755_0 ? _T_536_0_23 : _GEN_74;
  assign _GEN_76 = 5'h18 == _T_755_0 ? _T_536_0_24 : _GEN_75;
  assign _GEN_77 = 5'h19 == _T_755_0 ? _T_536_0_25 : _GEN_76;
  assign _GEN_78 = 5'h1a == _T_755_0 ? _T_536_0_26 : _GEN_77;
  assign _GEN_79 = 5'h1b == _T_755_0 ? _T_536_0_27 : _GEN_78;
  assign _GEN_80 = 5'h1c == _T_755_0 ? _T_536_0_28 : _GEN_79;
  assign _GEN_81 = 5'h1d == _T_755_0 ? _T_536_0_29 : _GEN_80;
  assign _GEN_82 = 5'h1e == _T_755_0 ? _T_536_0_30 : _GEN_81;
  assign _GEN_83 = 5'h1f == _T_755_0 ? _T_536_0_31 : _GEN_82;
  assign _T_4192 = _T_4144 ? _T_776_0 : 1'h0;
  assign _T_4197 = _T_4195 != 1'h1;
  assign _T_4199 = _T_4195 + 1'h1;
  assign _T_4200 = _T_4199[0:0];
  assign _GEN_84 = _T_4197 ? _T_4200 : _T_4195;
  assign _T_4208 = io_inputMemAddrReadys_1 | _T_309_0;
  assign _T_4209 = _T_4195 & _T_4208;
  assign _T_4211 = _T_4203 == 1'h0;
  assign _T_4216 = _T_245 + 1'h1;
  assign _T_4217 = _T_4216[0:0];
  assign _T_4218 = _T_245 ? 1'h1 : _T_4217;
  assign _T_4222 = _T_4203 + 1'h1;
  assign _T_4223 = _T_4222[0:0];
  assign _GEN_85 = _T_4211 ? _T_4218 : _T_245;
  assign _GEN_86 = _T_4211 ? 1'h0 : _GEN_84;
  assign _GEN_87 = _T_4211 ? 1'h0 : _T_4223;
  assign _GEN_88 = _T_4209 ? _GEN_85 : _T_245;
  assign _GEN_89 = _T_4209 ? _GEN_86 : _GEN_84;
  assign _GEN_90 = _T_4209 ? _GEN_87 : _T_4203;
  assign _T_4231 = _T_309_0 == 1'h0;
  assign _T_4232 = _T_4195 & _T_4231;
  assign _T_4237 = _T_4235 != 1'h1;
  assign _T_4239 = _T_4235 + 1'h1;
  assign _T_4240 = _T_4239[0:0];
  assign _GEN_91 = _T_4237 ? _T_4240 : _T_4235;
  assign _T_4570 = _T_4564 == 1'h0;
  assign _T_4571 = _T_4235 & _T_4570;
  assign _T_4572 = io_inputMemBlockReadys_1 & io_inputMemBlockValids_1;
  assign _T_4575 = _T_4572 | _T_315_0;
  assign _T_4576 = _T_4571 & _T_4575;
  assign _T_4680 = io_inputMemBlocks_1[15:0];
  assign _T_4784 = io_inputMemBlocks_1[31:16];
  assign _T_4888 = io_inputMemBlocks_1[47:32];
  assign _T_4992 = io_inputMemBlocks_1[63:48];
  assign _T_5096 = io_inputMemBlocks_1[79:64];
  assign _T_5200 = io_inputMemBlocks_1[95:80];
  assign _T_5304 = io_inputMemBlocks_1[111:96];
  assign _T_5408 = io_inputMemBlocks_1[127:112];
  assign _T_5512 = io_inputMemBlocks_1[143:128];
  assign _T_5616 = io_inputMemBlocks_1[159:144];
  assign _T_5720 = io_inputMemBlocks_1[175:160];
  assign _T_5824 = io_inputMemBlocks_1[191:176];
  assign _T_5928 = io_inputMemBlocks_1[207:192];
  assign _T_6032 = io_inputMemBlocks_1[223:208];
  assign _T_6136 = io_inputMemBlocks_1[239:224];
  assign _T_6240 = io_inputMemBlocks_1[255:240];
  assign _T_6344 = io_inputMemBlocks_1[271:256];
  assign _T_6448 = io_inputMemBlocks_1[287:272];
  assign _T_6552 = io_inputMemBlocks_1[303:288];
  assign _T_6656 = io_inputMemBlocks_1[319:304];
  assign _T_6760 = io_inputMemBlocks_1[335:320];
  assign _T_6864 = io_inputMemBlocks_1[351:336];
  assign _T_6968 = io_inputMemBlocks_1[367:352];
  assign _T_7072 = io_inputMemBlocks_1[383:368];
  assign _T_7176 = io_inputMemBlocks_1[399:384];
  assign _T_7280 = io_inputMemBlocks_1[415:400];
  assign _T_7384 = io_inputMemBlocks_1[431:416];
  assign _T_7488 = io_inputMemBlocks_1[447:432];
  assign _T_7592 = io_inputMemBlocks_1[463:448];
  assign _T_7696 = io_inputMemBlocks_1[479:464];
  assign _T_7800 = io_inputMemBlocks_1[495:480];
  assign _T_7904 = io_inputMemBlocks_1[511:496];
  assign _T_7912 = _T_315_0 == 1'h0;
  assign _T_7914 = _T_4564 + 1'h1;
  assign _T_7915 = _T_7914[0:0];
  assign _GEN_92 = _T_4576 ? _T_4680 : _T_4314_0_0;
  assign _GEN_93 = _T_4576 ? _T_4784 : _T_4314_0_1;
  assign _GEN_94 = _T_4576 ? _T_4888 : _T_4314_0_2;
  assign _GEN_95 = _T_4576 ? _T_4992 : _T_4314_0_3;
  assign _GEN_96 = _T_4576 ? _T_5096 : _T_4314_0_4;
  assign _GEN_97 = _T_4576 ? _T_5200 : _T_4314_0_5;
  assign _GEN_98 = _T_4576 ? _T_5304 : _T_4314_0_6;
  assign _GEN_99 = _T_4576 ? _T_5408 : _T_4314_0_7;
  assign _GEN_100 = _T_4576 ? _T_5512 : _T_4314_0_8;
  assign _GEN_101 = _T_4576 ? _T_5616 : _T_4314_0_9;
  assign _GEN_102 = _T_4576 ? _T_5720 : _T_4314_0_10;
  assign _GEN_103 = _T_4576 ? _T_5824 : _T_4314_0_11;
  assign _GEN_104 = _T_4576 ? _T_5928 : _T_4314_0_12;
  assign _GEN_105 = _T_4576 ? _T_6032 : _T_4314_0_13;
  assign _GEN_106 = _T_4576 ? _T_6136 : _T_4314_0_14;
  assign _GEN_107 = _T_4576 ? _T_6240 : _T_4314_0_15;
  assign _GEN_108 = _T_4576 ? _T_6344 : _T_4314_0_16;
  assign _GEN_109 = _T_4576 ? _T_6448 : _T_4314_0_17;
  assign _GEN_110 = _T_4576 ? _T_6552 : _T_4314_0_18;
  assign _GEN_111 = _T_4576 ? _T_6656 : _T_4314_0_19;
  assign _GEN_112 = _T_4576 ? _T_6760 : _T_4314_0_20;
  assign _GEN_113 = _T_4576 ? _T_6864 : _T_4314_0_21;
  assign _GEN_114 = _T_4576 ? _T_6968 : _T_4314_0_22;
  assign _GEN_115 = _T_4576 ? _T_7072 : _T_4314_0_23;
  assign _GEN_116 = _T_4576 ? _T_7176 : _T_4314_0_24;
  assign _GEN_117 = _T_4576 ? _T_7280 : _T_4314_0_25;
  assign _GEN_118 = _T_4576 ? _T_7384 : _T_4314_0_26;
  assign _GEN_119 = _T_4576 ? _T_7488 : _T_4314_0_27;
  assign _GEN_120 = _T_4576 ? _T_7592 : _T_4314_0_28;
  assign _GEN_121 = _T_4576 ? _T_7696 : _T_4314_0_29;
  assign _GEN_122 = _T_4576 ? _T_7800 : _T_4314_0_30;
  assign _GEN_123 = _T_4576 ? _T_7904 : _T_4314_0_31;
  assign _GEN_124 = _T_4576 ? _T_7912 : _T_4554_0;
  assign _GEN_125 = _T_4576 ? _T_7915 : _T_4564;
  assign _T_7919 = _T_4554_0 == 1'h0;
  assign _T_7920 = _T_4564 & _T_7919;
  assign _T_7925 = _T_248 + 1'h1;
  assign _T_7926 = _T_7925[0:0];
  assign _T_7927 = _T_248 ? 1'h1 : _T_7926;
  assign _GEN_126 = _T_7920 ? _T_7927 : _T_248;
  assign _GEN_127 = _T_7920 ? 1'h0 : _GEN_91;
  assign _GEN_128 = _T_7920 ? 1'h0 : _GEN_125;
  assign _T_7931 = {_T_248,_T_4564};
  assign _T_7936 = _T_4533_0 == 5'h1f;
  assign _T_7940 = _T_4533_0 + 5'h1;
  assign _T_7941 = _T_7940[4:0];
  assign _GEN_129 = _T_7936 ? 1'h0 : _GEN_124;
  assign _GEN_130 = _T_7936 ? 5'h0 : _T_7941;
  assign _GEN_131 = _T_4554_0 ? _GEN_129 : _GEN_124;
  assign _GEN_132 = _T_4554_0 ? _GEN_130 : _T_4533_0;
  assign _T_7951 = _T_4571 & _T_303_0;
  assign _T_7956 = _T_7951 & _T_7912;
  assign _T_7961 = _T_4211 & io_inputMemAddrReadys_1;
  assign _T_7962 = _T_7961 & io_inputMemAddrValids_1;
  assign _T_7964 = _T_245 ? _T_7962 : 1'h0;
  assign _GEN_133 = 5'h1 == _T_4533_0 ? _T_4314_0_1 : _T_4314_0_0;
  assign _GEN_134 = 5'h2 == _T_4533_0 ? _T_4314_0_2 : _GEN_133;
  assign _GEN_135 = 5'h3 == _T_4533_0 ? _T_4314_0_3 : _GEN_134;
  assign _GEN_136 = 5'h4 == _T_4533_0 ? _T_4314_0_4 : _GEN_135;
  assign _GEN_137 = 5'h5 == _T_4533_0 ? _T_4314_0_5 : _GEN_136;
  assign _GEN_138 = 5'h6 == _T_4533_0 ? _T_4314_0_6 : _GEN_137;
  assign _GEN_139 = 5'h7 == _T_4533_0 ? _T_4314_0_7 : _GEN_138;
  assign _GEN_140 = 5'h8 == _T_4533_0 ? _T_4314_0_8 : _GEN_139;
  assign _GEN_141 = 5'h9 == _T_4533_0 ? _T_4314_0_9 : _GEN_140;
  assign _GEN_142 = 5'ha == _T_4533_0 ? _T_4314_0_10 : _GEN_141;
  assign _GEN_143 = 5'hb == _T_4533_0 ? _T_4314_0_11 : _GEN_142;
  assign _GEN_144 = 5'hc == _T_4533_0 ? _T_4314_0_12 : _GEN_143;
  assign _GEN_145 = 5'hd == _T_4533_0 ? _T_4314_0_13 : _GEN_144;
  assign _GEN_146 = 5'he == _T_4533_0 ? _T_4314_0_14 : _GEN_145;
  assign _GEN_147 = 5'hf == _T_4533_0 ? _T_4314_0_15 : _GEN_146;
  assign _GEN_148 = 5'h10 == _T_4533_0 ? _T_4314_0_16 : _GEN_147;
  assign _GEN_149 = 5'h11 == _T_4533_0 ? _T_4314_0_17 : _GEN_148;
  assign _GEN_150 = 5'h12 == _T_4533_0 ? _T_4314_0_18 : _GEN_149;
  assign _GEN_151 = 5'h13 == _T_4533_0 ? _T_4314_0_19 : _GEN_150;
  assign _GEN_152 = 5'h14 == _T_4533_0 ? _T_4314_0_20 : _GEN_151;
  assign _GEN_153 = 5'h15 == _T_4533_0 ? _T_4314_0_21 : _GEN_152;
  assign _GEN_154 = 5'h16 == _T_4533_0 ? _T_4314_0_22 : _GEN_153;
  assign _GEN_155 = 5'h17 == _T_4533_0 ? _T_4314_0_23 : _GEN_154;
  assign _GEN_156 = 5'h18 == _T_4533_0 ? _T_4314_0_24 : _GEN_155;
  assign _GEN_157 = 5'h19 == _T_4533_0 ? _T_4314_0_25 : _GEN_156;
  assign _GEN_158 = 5'h1a == _T_4533_0 ? _T_4314_0_26 : _GEN_157;
  assign _GEN_159 = 5'h1b == _T_4533_0 ? _T_4314_0_27 : _GEN_158;
  assign _GEN_160 = 5'h1c == _T_4533_0 ? _T_4314_0_28 : _GEN_159;
  assign _GEN_161 = 5'h1d == _T_4533_0 ? _T_4314_0_29 : _GEN_160;
  assign _GEN_162 = 5'h1e == _T_4533_0 ? _T_4314_0_30 : _GEN_161;
  assign _GEN_163 = 5'h1f == _T_4533_0 ? _T_4314_0_31 : _GEN_162;
  assign _T_7970 = _T_248 ? _T_4554_0 : 1'h0;
  assign _T_7975 = _T_7973 != 1'h1;
  assign _T_7977 = _T_7973 + 1'h1;
  assign _T_7978 = _T_7977[0:0];
  assign _GEN_164 = _T_7975 ? _T_7978 : _T_7973;
  assign _T_8319 = _T_8315 == 1'h0;
  assign _T_8320 = _T_7973 & _T_8319;
  assign _GEN_165 = _T_8320 ? 1'h1 : _T_8315;
  assign _T_8324 = _T_7973 & _T_345_0;
  assign _T_8326 = _T_357_0 == 5'h1f;
  assign _T_8327 = _T_8324 & _T_8326;
  assign _GEN_166 = _T_8327 ? 1'h1 : _T_8299_0;
  assign _GEN_167 = 5'h0 == _T_357_0 ? _GEN_2 : _T_8080_0_0;
  assign _GEN_168 = 5'h1 == _T_357_0 ? _GEN_2 : _T_8080_0_1;
  assign _GEN_169 = 5'h2 == _T_357_0 ? _GEN_2 : _T_8080_0_2;
  assign _GEN_170 = 5'h3 == _T_357_0 ? _GEN_2 : _T_8080_0_3;
  assign _GEN_171 = 5'h4 == _T_357_0 ? _GEN_2 : _T_8080_0_4;
  assign _GEN_172 = 5'h5 == _T_357_0 ? _GEN_2 : _T_8080_0_5;
  assign _GEN_173 = 5'h6 == _T_357_0 ? _GEN_2 : _T_8080_0_6;
  assign _GEN_174 = 5'h7 == _T_357_0 ? _GEN_2 : _T_8080_0_7;
  assign _GEN_175 = 5'h8 == _T_357_0 ? _GEN_2 : _T_8080_0_8;
  assign _GEN_176 = 5'h9 == _T_357_0 ? _GEN_2 : _T_8080_0_9;
  assign _GEN_177 = 5'ha == _T_357_0 ? _GEN_2 : _T_8080_0_10;
  assign _GEN_178 = 5'hb == _T_357_0 ? _GEN_2 : _T_8080_0_11;
  assign _GEN_179 = 5'hc == _T_357_0 ? _GEN_2 : _T_8080_0_12;
  assign _GEN_180 = 5'hd == _T_357_0 ? _GEN_2 : _T_8080_0_13;
  assign _GEN_181 = 5'he == _T_357_0 ? _GEN_2 : _T_8080_0_14;
  assign _GEN_182 = 5'hf == _T_357_0 ? _GEN_2 : _T_8080_0_15;
  assign _GEN_183 = 5'h10 == _T_357_0 ? _GEN_2 : _T_8080_0_16;
  assign _GEN_184 = 5'h11 == _T_357_0 ? _GEN_2 : _T_8080_0_17;
  assign _GEN_185 = 5'h12 == _T_357_0 ? _GEN_2 : _T_8080_0_18;
  assign _GEN_186 = 5'h13 == _T_357_0 ? _GEN_2 : _T_8080_0_19;
  assign _GEN_187 = 5'h14 == _T_357_0 ? _GEN_2 : _T_8080_0_20;
  assign _GEN_188 = 5'h15 == _T_357_0 ? _GEN_2 : _T_8080_0_21;
  assign _GEN_189 = 5'h16 == _T_357_0 ? _GEN_2 : _T_8080_0_22;
  assign _GEN_190 = 5'h17 == _T_357_0 ? _GEN_2 : _T_8080_0_23;
  assign _GEN_191 = 5'h18 == _T_357_0 ? _GEN_2 : _T_8080_0_24;
  assign _GEN_192 = 5'h19 == _T_357_0 ? _GEN_2 : _T_8080_0_25;
  assign _GEN_193 = 5'h1a == _T_357_0 ? _GEN_2 : _T_8080_0_26;
  assign _GEN_194 = 5'h1b == _T_357_0 ? _GEN_2 : _T_8080_0_27;
  assign _GEN_195 = 5'h1c == _T_357_0 ? _GEN_2 : _T_8080_0_28;
  assign _GEN_196 = 5'h1d == _T_357_0 ? _GEN_2 : _T_8080_0_29;
  assign _GEN_197 = 5'h1e == _T_357_0 ? _GEN_2 : _T_8080_0_30;
  assign _GEN_198 = 5'h1f == _T_357_0 ? _GEN_2 : _T_8080_0_31;
  assign _GEN_199 = _T_345_0 ? _GEN_167 : _T_8080_0_0;
  assign _GEN_200 = _T_345_0 ? _GEN_168 : _T_8080_0_1;
  assign _GEN_201 = _T_345_0 ? _GEN_169 : _T_8080_0_2;
  assign _GEN_202 = _T_345_0 ? _GEN_170 : _T_8080_0_3;
  assign _GEN_203 = _T_345_0 ? _GEN_171 : _T_8080_0_4;
  assign _GEN_204 = _T_345_0 ? _GEN_172 : _T_8080_0_5;
  assign _GEN_205 = _T_345_0 ? _GEN_173 : _T_8080_0_6;
  assign _GEN_206 = _T_345_0 ? _GEN_174 : _T_8080_0_7;
  assign _GEN_207 = _T_345_0 ? _GEN_175 : _T_8080_0_8;
  assign _GEN_208 = _T_345_0 ? _GEN_176 : _T_8080_0_9;
  assign _GEN_209 = _T_345_0 ? _GEN_177 : _T_8080_0_10;
  assign _GEN_210 = _T_345_0 ? _GEN_178 : _T_8080_0_11;
  assign _GEN_211 = _T_345_0 ? _GEN_179 : _T_8080_0_12;
  assign _GEN_212 = _T_345_0 ? _GEN_180 : _T_8080_0_13;
  assign _GEN_213 = _T_345_0 ? _GEN_181 : _T_8080_0_14;
  assign _GEN_214 = _T_345_0 ? _GEN_182 : _T_8080_0_15;
  assign _GEN_215 = _T_345_0 ? _GEN_183 : _T_8080_0_16;
  assign _GEN_216 = _T_345_0 ? _GEN_184 : _T_8080_0_17;
  assign _GEN_217 = _T_345_0 ? _GEN_185 : _T_8080_0_18;
  assign _GEN_218 = _T_345_0 ? _GEN_186 : _T_8080_0_19;
  assign _GEN_219 = _T_345_0 ? _GEN_187 : _T_8080_0_20;
  assign _GEN_220 = _T_345_0 ? _GEN_188 : _T_8080_0_21;
  assign _GEN_221 = _T_345_0 ? _GEN_189 : _T_8080_0_22;
  assign _GEN_222 = _T_345_0 ? _GEN_190 : _T_8080_0_23;
  assign _GEN_223 = _T_345_0 ? _GEN_191 : _T_8080_0_24;
  assign _GEN_224 = _T_345_0 ? _GEN_192 : _T_8080_0_25;
  assign _GEN_225 = _T_345_0 ? _GEN_193 : _T_8080_0_26;
  assign _GEN_226 = _T_345_0 ? _GEN_194 : _T_8080_0_27;
  assign _GEN_227 = _T_345_0 ? _GEN_195 : _T_8080_0_28;
  assign _GEN_228 = _T_345_0 ? _GEN_196 : _T_8080_0_29;
  assign _GEN_229 = _T_345_0 ? _GEN_197 : _T_8080_0_30;
  assign _GEN_230 = _T_345_0 ? _GEN_198 : _T_8080_0_31;
  assign _T_8333 = _T_7973 & _T_339_0;
  assign _T_8335 = _T_7992_0 == 1'h0;
  assign _T_8336 = _T_8333 & _T_8335;
  assign _T_8342 = _T_8336 & _T_8319;
  assign _GEN_231 = _T_8342 ? 1'h1 : _T_7992_0;
  assign _GEN_232 = _T_8342 ? _T_333_0 : _T_8003_0;
  assign _T_8351 = _T_8312 == 1'h0;
  assign _T_8352 = _T_7992_0 & _T_8351;
  assign _T_8456 = {_T_8080_0_1,_T_8080_0_0};
  assign _T_8457 = {_T_8080_0_3,_T_8080_0_2};
  assign _T_8458 = {_T_8457,_T_8456};
  assign _T_8459 = {_T_8080_0_5,_T_8080_0_4};
  assign _T_8460 = {_T_8080_0_7,_T_8080_0_6};
  assign _T_8461 = {_T_8460,_T_8459};
  assign _T_8462 = {_T_8461,_T_8458};
  assign _T_8463 = {_T_8080_0_9,_T_8080_0_8};
  assign _T_8464 = {_T_8080_0_11,_T_8080_0_10};
  assign _T_8465 = {_T_8464,_T_8463};
  assign _T_8466 = {_T_8080_0_13,_T_8080_0_12};
  assign _T_8467 = {_T_8080_0_15,_T_8080_0_14};
  assign _T_8468 = {_T_8467,_T_8466};
  assign _T_8469 = {_T_8468,_T_8465};
  assign _T_8470 = {_T_8469,_T_8462};
  assign _T_8471 = {_T_8080_0_17,_T_8080_0_16};
  assign _T_8472 = {_T_8080_0_19,_T_8080_0_18};
  assign _T_8473 = {_T_8472,_T_8471};
  assign _T_8474 = {_T_8080_0_21,_T_8080_0_20};
  assign _T_8475 = {_T_8080_0_23,_T_8080_0_22};
  assign _T_8476 = {_T_8475,_T_8474};
  assign _T_8477 = {_T_8476,_T_8473};
  assign _T_8478 = {_T_8080_0_25,_T_8080_0_24};
  assign _T_8479 = {_T_8080_0_27,_T_8080_0_26};
  assign _T_8480 = {_T_8479,_T_8478};
  assign _T_8481 = {_T_8080_0_29,_T_8080_0_28};
  assign _T_8482 = {_T_8080_0_31,_T_8080_0_30};
  assign _T_8483 = {_T_8482,_T_8481};
  assign _T_8484 = {_T_8483,_T_8480};
  assign _T_8485 = {_T_8484,_T_8477};
  assign _T_8486 = {_T_8485,_T_8470};
  assign _T_8491 = _T_8299_0 & _T_8312;
  assign _T_8498 = _T_7973 & _T_363_0;
  assign _T_8501 = io_outputMemAddrValids_0 & io_outputMemAddrReadys_0;
  assign _T_8502 = _T_8493 | _T_8501;
  assign _T_8509 = _T_8315 & _T_8335;
  assign _T_8510 = _T_8502 | _T_8509;
  assign _T_8511 = _T_8351 & _T_8510;
  assign _GEN_233 = _T_8511 ? 1'h1 : _T_8312;
  assign _T_8513 = io_outputMemBlockValids_0 & io_outputMemBlockReadys_0;
  assign _T_8514 = _T_8493 | _T_8513;
  assign _T_8521 = _T_8514 | _T_8335;
  assign _T_8522 = _T_8312 & _T_8521;
  assign _T_8525 = _T_8309 == 1'h0;
  assign _T_8527 = _T_251 == 1'h0;
  assign _T_8530 = _T_251 + 1'h1;
  assign _T_8531 = _T_8530[0:0];
  assign _T_8532 = _T_8527 ? 1'h0 : _T_8531;
  assign _T_8539 = _T_8309 + 1'h1;
  assign _T_8540 = _T_8539[0:0];
  assign _GEN_234 = _T_8525 ? _T_8532 : _T_251;
  assign _GEN_235 = _T_8525 ? 1'h0 : _GEN_164;
  assign _GEN_236 = _T_8525 ? 1'h0 : _T_8540;
  assign _GEN_237 = _T_8525 ? 1'h0 : _GEN_165;
  assign _GEN_238 = _T_8525 ? 1'h0 : _GEN_231;
  assign _GEN_239 = _T_8525 ? 1'h0 : _GEN_166;
  assign _GEN_240 = _T_8522 ? 1'h0 : _GEN_233;
  assign _GEN_241 = _T_8522 ? _GEN_234 : _T_251;
  assign _GEN_242 = _T_8522 ? _GEN_235 : _GEN_164;
  assign _GEN_243 = _T_8522 ? _GEN_236 : _T_8309;
  assign _GEN_244 = _T_8522 ? _GEN_237 : _GEN_165;
  assign _GEN_245 = _T_8522 ? _GEN_238 : _GEN_231;
  assign _GEN_246 = _T_8522 ? _GEN_239 : _GEN_166;
  assign _T_8556 = _T_8527 ? _T_8342 : 1'h0;
  assign _T_8561 = _T_8525 & io_outputMemBlockValids_0;
  assign _T_8562 = _T_8561 & io_outputMemBlockReadys_0;
  assign _T_8564 = _T_8527 ? _T_8562 : 1'h0;
  assign _T_8565 = io_outputMemBlockReadys_0 & io_outputMemBlockValids_0;
  assign _T_8566 = {_T_251,_T_8309};
  assign _T_8574 = _T_8572 != 1'h1;
  assign _T_8576 = _T_8572 + 1'h1;
  assign _T_8577 = _T_8576[0:0];
  assign _GEN_247 = _T_8574 ? _T_8577 : _T_8572;
  assign _T_8918 = _T_8914 == 1'h0;
  assign _T_8919 = _T_8572 & _T_8918;
  assign _GEN_248 = _T_8919 ? 1'h1 : _T_8914;
  assign _T_8923 = _T_8572 & _T_393_0;
  assign _T_8925 = _T_405_0 == 5'h1f;
  assign _T_8926 = _T_8923 & _T_8925;
  assign _GEN_249 = _T_8926 ? 1'h1 : _T_8898_0;
  assign _GEN_250 = 5'h0 == _T_405_0 ? _GEN_3 : _T_8679_0_0;
  assign _GEN_251 = 5'h1 == _T_405_0 ? _GEN_3 : _T_8679_0_1;
  assign _GEN_252 = 5'h2 == _T_405_0 ? _GEN_3 : _T_8679_0_2;
  assign _GEN_253 = 5'h3 == _T_405_0 ? _GEN_3 : _T_8679_0_3;
  assign _GEN_254 = 5'h4 == _T_405_0 ? _GEN_3 : _T_8679_0_4;
  assign _GEN_255 = 5'h5 == _T_405_0 ? _GEN_3 : _T_8679_0_5;
  assign _GEN_256 = 5'h6 == _T_405_0 ? _GEN_3 : _T_8679_0_6;
  assign _GEN_257 = 5'h7 == _T_405_0 ? _GEN_3 : _T_8679_0_7;
  assign _GEN_258 = 5'h8 == _T_405_0 ? _GEN_3 : _T_8679_0_8;
  assign _GEN_259 = 5'h9 == _T_405_0 ? _GEN_3 : _T_8679_0_9;
  assign _GEN_260 = 5'ha == _T_405_0 ? _GEN_3 : _T_8679_0_10;
  assign _GEN_261 = 5'hb == _T_405_0 ? _GEN_3 : _T_8679_0_11;
  assign _GEN_262 = 5'hc == _T_405_0 ? _GEN_3 : _T_8679_0_12;
  assign _GEN_263 = 5'hd == _T_405_0 ? _GEN_3 : _T_8679_0_13;
  assign _GEN_264 = 5'he == _T_405_0 ? _GEN_3 : _T_8679_0_14;
  assign _GEN_265 = 5'hf == _T_405_0 ? _GEN_3 : _T_8679_0_15;
  assign _GEN_266 = 5'h10 == _T_405_0 ? _GEN_3 : _T_8679_0_16;
  assign _GEN_267 = 5'h11 == _T_405_0 ? _GEN_3 : _T_8679_0_17;
  assign _GEN_268 = 5'h12 == _T_405_0 ? _GEN_3 : _T_8679_0_18;
  assign _GEN_269 = 5'h13 == _T_405_0 ? _GEN_3 : _T_8679_0_19;
  assign _GEN_270 = 5'h14 == _T_405_0 ? _GEN_3 : _T_8679_0_20;
  assign _GEN_271 = 5'h15 == _T_405_0 ? _GEN_3 : _T_8679_0_21;
  assign _GEN_272 = 5'h16 == _T_405_0 ? _GEN_3 : _T_8679_0_22;
  assign _GEN_273 = 5'h17 == _T_405_0 ? _GEN_3 : _T_8679_0_23;
  assign _GEN_274 = 5'h18 == _T_405_0 ? _GEN_3 : _T_8679_0_24;
  assign _GEN_275 = 5'h19 == _T_405_0 ? _GEN_3 : _T_8679_0_25;
  assign _GEN_276 = 5'h1a == _T_405_0 ? _GEN_3 : _T_8679_0_26;
  assign _GEN_277 = 5'h1b == _T_405_0 ? _GEN_3 : _T_8679_0_27;
  assign _GEN_278 = 5'h1c == _T_405_0 ? _GEN_3 : _T_8679_0_28;
  assign _GEN_279 = 5'h1d == _T_405_0 ? _GEN_3 : _T_8679_0_29;
  assign _GEN_280 = 5'h1e == _T_405_0 ? _GEN_3 : _T_8679_0_30;
  assign _GEN_281 = 5'h1f == _T_405_0 ? _GEN_3 : _T_8679_0_31;
  assign _GEN_282 = _T_393_0 ? _GEN_250 : _T_8679_0_0;
  assign _GEN_283 = _T_393_0 ? _GEN_251 : _T_8679_0_1;
  assign _GEN_284 = _T_393_0 ? _GEN_252 : _T_8679_0_2;
  assign _GEN_285 = _T_393_0 ? _GEN_253 : _T_8679_0_3;
  assign _GEN_286 = _T_393_0 ? _GEN_254 : _T_8679_0_4;
  assign _GEN_287 = _T_393_0 ? _GEN_255 : _T_8679_0_5;
  assign _GEN_288 = _T_393_0 ? _GEN_256 : _T_8679_0_6;
  assign _GEN_289 = _T_393_0 ? _GEN_257 : _T_8679_0_7;
  assign _GEN_290 = _T_393_0 ? _GEN_258 : _T_8679_0_8;
  assign _GEN_291 = _T_393_0 ? _GEN_259 : _T_8679_0_9;
  assign _GEN_292 = _T_393_0 ? _GEN_260 : _T_8679_0_10;
  assign _GEN_293 = _T_393_0 ? _GEN_261 : _T_8679_0_11;
  assign _GEN_294 = _T_393_0 ? _GEN_262 : _T_8679_0_12;
  assign _GEN_295 = _T_393_0 ? _GEN_263 : _T_8679_0_13;
  assign _GEN_296 = _T_393_0 ? _GEN_264 : _T_8679_0_14;
  assign _GEN_297 = _T_393_0 ? _GEN_265 : _T_8679_0_15;
  assign _GEN_298 = _T_393_0 ? _GEN_266 : _T_8679_0_16;
  assign _GEN_299 = _T_393_0 ? _GEN_267 : _T_8679_0_17;
  assign _GEN_300 = _T_393_0 ? _GEN_268 : _T_8679_0_18;
  assign _GEN_301 = _T_393_0 ? _GEN_269 : _T_8679_0_19;
  assign _GEN_302 = _T_393_0 ? _GEN_270 : _T_8679_0_20;
  assign _GEN_303 = _T_393_0 ? _GEN_271 : _T_8679_0_21;
  assign _GEN_304 = _T_393_0 ? _GEN_272 : _T_8679_0_22;
  assign _GEN_305 = _T_393_0 ? _GEN_273 : _T_8679_0_23;
  assign _GEN_306 = _T_393_0 ? _GEN_274 : _T_8679_0_24;
  assign _GEN_307 = _T_393_0 ? _GEN_275 : _T_8679_0_25;
  assign _GEN_308 = _T_393_0 ? _GEN_276 : _T_8679_0_26;
  assign _GEN_309 = _T_393_0 ? _GEN_277 : _T_8679_0_27;
  assign _GEN_310 = _T_393_0 ? _GEN_278 : _T_8679_0_28;
  assign _GEN_311 = _T_393_0 ? _GEN_279 : _T_8679_0_29;
  assign _GEN_312 = _T_393_0 ? _GEN_280 : _T_8679_0_30;
  assign _GEN_313 = _T_393_0 ? _GEN_281 : _T_8679_0_31;
  assign _T_8932 = _T_8572 & _T_387_0;
  assign _T_8934 = _T_8591_0 == 1'h0;
  assign _T_8935 = _T_8932 & _T_8934;
  assign _T_8941 = _T_8935 & _T_8918;
  assign _GEN_314 = _T_8941 ? 1'h1 : _T_8591_0;
  assign _GEN_315 = _T_8941 ? _T_381_0 : _T_8602_0;
  assign _T_8950 = _T_8911 == 1'h0;
  assign _T_8951 = _T_8591_0 & _T_8950;
  assign _T_9055 = {_T_8679_0_1,_T_8679_0_0};
  assign _T_9056 = {_T_8679_0_3,_T_8679_0_2};
  assign _T_9057 = {_T_9056,_T_9055};
  assign _T_9058 = {_T_8679_0_5,_T_8679_0_4};
  assign _T_9059 = {_T_8679_0_7,_T_8679_0_6};
  assign _T_9060 = {_T_9059,_T_9058};
  assign _T_9061 = {_T_9060,_T_9057};
  assign _T_9062 = {_T_8679_0_9,_T_8679_0_8};
  assign _T_9063 = {_T_8679_0_11,_T_8679_0_10};
  assign _T_9064 = {_T_9063,_T_9062};
  assign _T_9065 = {_T_8679_0_13,_T_8679_0_12};
  assign _T_9066 = {_T_8679_0_15,_T_8679_0_14};
  assign _T_9067 = {_T_9066,_T_9065};
  assign _T_9068 = {_T_9067,_T_9064};
  assign _T_9069 = {_T_9068,_T_9061};
  assign _T_9070 = {_T_8679_0_17,_T_8679_0_16};
  assign _T_9071 = {_T_8679_0_19,_T_8679_0_18};
  assign _T_9072 = {_T_9071,_T_9070};
  assign _T_9073 = {_T_8679_0_21,_T_8679_0_20};
  assign _T_9074 = {_T_8679_0_23,_T_8679_0_22};
  assign _T_9075 = {_T_9074,_T_9073};
  assign _T_9076 = {_T_9075,_T_9072};
  assign _T_9077 = {_T_8679_0_25,_T_8679_0_24};
  assign _T_9078 = {_T_8679_0_27,_T_8679_0_26};
  assign _T_9079 = {_T_9078,_T_9077};
  assign _T_9080 = {_T_8679_0_29,_T_8679_0_28};
  assign _T_9081 = {_T_8679_0_31,_T_8679_0_30};
  assign _T_9082 = {_T_9081,_T_9080};
  assign _T_9083 = {_T_9082,_T_9079};
  assign _T_9084 = {_T_9083,_T_9076};
  assign _T_9085 = {_T_9084,_T_9069};
  assign _T_9090 = _T_8898_0 & _T_8911;
  assign _T_9097 = _T_8572 & _T_411_0;
  assign _T_9100 = io_outputMemAddrValids_1 & io_outputMemAddrReadys_1;
  assign _T_9101 = _T_9092 | _T_9100;
  assign _T_9108 = _T_8914 & _T_8934;
  assign _T_9109 = _T_9101 | _T_9108;
  assign _T_9110 = _T_8950 & _T_9109;
  assign _GEN_316 = _T_9110 ? 1'h1 : _T_8911;
  assign _T_9112 = io_outputMemBlockValids_1 & io_outputMemBlockReadys_1;
  assign _T_9113 = _T_9092 | _T_9112;
  assign _T_9120 = _T_9113 | _T_8934;
  assign _T_9121 = _T_8911 & _T_9120;
  assign _T_9124 = _T_8908 == 1'h0;
  assign _T_9129 = _T_254 + 1'h1;
  assign _T_9130 = _T_9129[0:0];
  assign _T_9131 = _T_254 ? 1'h1 : _T_9130;
  assign _T_9138 = _T_8908 + 1'h1;
  assign _T_9139 = _T_9138[0:0];
  assign _GEN_317 = _T_9124 ? _T_9131 : _T_254;
  assign _GEN_318 = _T_9124 ? 1'h0 : _GEN_247;
  assign _GEN_319 = _T_9124 ? 1'h0 : _T_9139;
  assign _GEN_320 = _T_9124 ? 1'h0 : _GEN_248;
  assign _GEN_321 = _T_9124 ? 1'h0 : _GEN_314;
  assign _GEN_322 = _T_9124 ? 1'h0 : _GEN_249;
  assign _GEN_323 = _T_9121 ? 1'h0 : _GEN_316;
  assign _GEN_324 = _T_9121 ? _GEN_317 : _T_254;
  assign _GEN_325 = _T_9121 ? _GEN_318 : _GEN_247;
  assign _GEN_326 = _T_9121 ? _GEN_319 : _T_8908;
  assign _GEN_327 = _T_9121 ? _GEN_320 : _GEN_248;
  assign _GEN_328 = _T_9121 ? _GEN_321 : _GEN_314;
  assign _GEN_329 = _T_9121 ? _GEN_322 : _GEN_249;
  assign _T_9155 = _T_254 ? _T_8941 : 1'h0;
  assign _T_9160 = _T_9124 & io_outputMemBlockValids_1;
  assign _T_9161 = _T_9160 & io_outputMemBlockReadys_1;
  assign _T_9163 = _T_254 ? _T_9161 : 1'h0;
  assign _T_9164 = io_outputMemBlockReadys_1 & io_outputMemBlockValids_1;
  assign _T_9165 = {_T_254,_T_8908};
  assign cumFinished = cores_0_outputFinished & cores_1_outputFinished;
  assign io_inputMemAddrs_0 = {{32'd0}, _T_265_0};
  assign io_inputMemAddrs_1 = {{32'd0}, _T_297_0};
  assign io_inputMemAddrValids_0 = _T_454;
  assign io_inputMemAddrValids_1 = _T_4232;
  assign io_inputMemBlockReadys_0 = _T_4178;
  assign io_inputMemBlockReadys_1 = _T_7956;
  assign io_outputMemAddrs_0 = {{32'd0}, _T_8003_0};
  assign io_outputMemAddrs_1 = {{32'd0}, _T_8602_0};
  assign io_outputMemAddrValids_0 = _T_8352;
  assign io_outputMemAddrValids_1 = _T_8951;
  assign io_outputMemBlocks_0 = _T_8486;
  assign io_outputMemBlocks_1 = _T_9085;
  assign io_outputMemBlockValids_0 = _T_8491;
  assign io_outputMemBlockValids_1 = _T_9090;
  assign io_finished = cumFinished;
  assign StreamingCore_io_inputMemAddrConsumed = cores_0_inputMemAddrConsumed;
  assign StreamingCore_io_inputMemBlock = cores_0_inputMemBlock;
  assign StreamingCore_io_inputMemIdx = cores_0_inputMemIdx;
  assign StreamingCore_io_inputMemBlockValid = cores_0_inputMemBlockValid;
  assign StreamingCore_io_outputMemAddrReady = cores_0_outputMemAddrReady;
  assign StreamingCore_io_outputMemBlockReady = cores_0_outputMemBlockReady;
  assign StreamingCore_clock = clock;
  assign StreamingCore_reset = reset;
  assign StreamingCore_1_io_inputMemAddrConsumed = cores_1_inputMemAddrConsumed;
  assign StreamingCore_1_io_inputMemBlock = cores_1_inputMemBlock;
  assign StreamingCore_1_io_inputMemIdx = cores_1_inputMemIdx;
  assign StreamingCore_1_io_inputMemBlockValid = cores_1_inputMemBlockValid;
  assign StreamingCore_1_io_outputMemAddrReady = cores_1_outputMemAddrReady;
  assign StreamingCore_1_io_outputMemBlockReady = cores_1_outputMemBlockReady;
  assign StreamingCore_1_clock = clock;
  assign StreamingCore_1_reset = reset;
  assign cores_0_inputMemAddr = StreamingCore_io_inputMemAddr;
  assign cores_0_inputMemAddrConsumed = _T_4186;
  assign cores_0_inputMemBlock = _GEN_0;
  assign cores_0_inputMemIdx = _T_755_0;
  assign cores_0_inputMemBlockValid = _T_4192;
  assign cores_0_inputMemBlockReady = StreamingCore_io_inputMemBlockReady;
  assign cores_0_outputMemAddr = StreamingCore_io_outputMemAddr;
  assign cores_0_outputMemAddrValid = StreamingCore_io_outputMemAddrValid;
  assign cores_0_outputMemAddrReady = _T_8556;
  assign cores_0_outputMemBlock = StreamingCore_io_outputMemBlock;
  assign cores_0_outputMemIdx = StreamingCore_io_outputMemIdx;
  assign cores_0_outputMemBlockValid = StreamingCore_io_outputMemBlockValid;
  assign cores_0_outputMemBlockReady = _T_8564;
  assign cores_0_inputAddrsIgnore = StreamingCore_io_inputAddrsIgnore;
  assign cores_0_inputBlocksFinished = StreamingCore_io_inputBlocksFinished;
  assign cores_0_outputFinished = StreamingCore_io_outputFinished;
  assign cores_1_inputMemAddr = StreamingCore_1_io_inputMemAddr;
  assign cores_1_inputMemAddrConsumed = _T_7964;
  assign cores_1_inputMemBlock = _GEN_1;
  assign cores_1_inputMemIdx = _T_4533_0;
  assign cores_1_inputMemBlockValid = _T_7970;
  assign cores_1_inputMemBlockReady = StreamingCore_1_io_inputMemBlockReady;
  assign cores_1_outputMemAddr = StreamingCore_1_io_outputMemAddr;
  assign cores_1_outputMemAddrValid = StreamingCore_1_io_outputMemAddrValid;
  assign cores_1_outputMemAddrReady = _T_9155;
  assign cores_1_outputMemBlock = StreamingCore_1_io_outputMemBlock;
  assign cores_1_outputMemIdx = StreamingCore_1_io_outputMemIdx;
  assign cores_1_outputMemBlockValid = StreamingCore_1_io_outputMemBlockValid;
  assign cores_1_outputMemBlockReady = _T_9163;
  assign cores_1_inputAddrsIgnore = StreamingCore_1_io_inputAddrsIgnore;
  assign cores_1_inputBlocksFinished = StreamingCore_1_io_inputBlocksFinished;
  assign cores_1_outputFinished = StreamingCore_1_io_outputFinished;
  assign _T_265_0 = _T_256;
  assign _T_271_0 = _T_258;
  assign _T_277_0 = _T_260;
  assign _T_283_0 = _T_262;
  assign _T_297_0 = _T_288;
  assign _T_303_0 = _T_290;
  assign _T_309_0 = _T_292;
  assign _T_315_0 = _T_294;
  assign _T_333_0 = _T_320;
  assign _T_339_0 = _T_322;
  assign _T_345_0 = _T_324;
  assign _T_351_0 = _T_326;
  assign _T_357_0 = _T_328;
  assign _T_363_0 = _T_330;
  assign _T_381_0 = _T_368;
  assign _T_387_0 = _T_370;
  assign _T_393_0 = _T_372;
  assign _T_399_0 = _T_374;
  assign _T_405_0 = _T_376;
  assign _T_411_0 = _T_378;
  assign _GEN_0 = _GEN_83;
  assign _GEN_1 = _GEN_163;
  assign _GEN_2 = _T_351_0;
  assign _T_8493 = _T_8498;
  assign _GEN_3 = _T_399_0;
  assign _T_9092 = _T_9097;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_239 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_242 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_245 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_248 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_251 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_254 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_256 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_258 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_260 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_262 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_288 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_290 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_292 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_294 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_320 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_322 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_324 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_326 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_328 = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_330 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_368 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_370 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_372 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_374 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_376 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_378 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_417 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_425 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_457 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_536_0_0 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_536_0_1 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_536_0_2 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_536_0_3 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_536_0_4 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_536_0_5 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_536_0_6 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_536_0_7 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_536_0_8 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_536_0_9 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_536_0_10 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_536_0_11 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_536_0_12 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_536_0_13 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_536_0_14 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_536_0_15 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_536_0_16 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_536_0_17 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_536_0_18 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_536_0_19 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_536_0_20 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_536_0_21 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_536_0_22 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_536_0_23 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_536_0_24 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_536_0_25 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_536_0_26 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_536_0_27 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_536_0_28 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_536_0_29 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_536_0_30 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_536_0_31 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_755_0 = _RAND_61[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_776_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_786 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_4195 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_4203 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_4235 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_4314_0_0 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_4314_0_1 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_4314_0_2 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_4314_0_3 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_4314_0_4 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_4314_0_5 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_4314_0_6 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_4314_0_7 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_4314_0_8 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_4314_0_9 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_4314_0_10 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_4314_0_11 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_4314_0_12 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_4314_0_13 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_4314_0_14 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_4314_0_15 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_4314_0_16 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_4314_0_17 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_4314_0_18 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_4314_0_19 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_4314_0_20 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_4314_0_21 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_4314_0_22 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_4314_0_23 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_4314_0_24 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_4314_0_25 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_4314_0_26 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_4314_0_27 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_4314_0_28 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_4314_0_29 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_4314_0_30 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_4314_0_31 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_4533_0 = _RAND_99[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_4554_0 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_4564 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_7973 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_7992_0 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_8003_0 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_8080_0_0 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_8080_0_1 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_8080_0_2 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_8080_0_3 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_8080_0_4 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_8080_0_5 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_8080_0_6 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_8080_0_7 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_8080_0_8 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_8080_0_9 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_8080_0_10 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_8080_0_11 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_8080_0_12 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_8080_0_13 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_8080_0_14 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_8080_0_15 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_8080_0_16 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_8080_0_17 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_8080_0_18 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_8080_0_19 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_8080_0_20 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_8080_0_21 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_8080_0_22 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_8080_0_23 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_8080_0_24 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_8080_0_25 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_8080_0_26 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_8080_0_27 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_8080_0_28 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_8080_0_29 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  _T_8080_0_30 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_8080_0_31 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  _T_8299_0 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  _T_8309 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  _T_8312 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  _T_8315 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  _T_8572 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  _T_8591_0 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  _T_8602_0 = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  _T_8679_0_0 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  _T_8679_0_1 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  _T_8679_0_2 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  _T_8679_0_3 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  _T_8679_0_4 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  _T_8679_0_5 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  _T_8679_0_6 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  _T_8679_0_7 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  _T_8679_0_8 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  _T_8679_0_9 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  _T_8679_0_10 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _T_8679_0_11 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  _T_8679_0_12 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _T_8679_0_13 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  _T_8679_0_14 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  _T_8679_0_15 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _T_8679_0_16 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  _T_8679_0_17 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  _T_8679_0_18 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  _T_8679_0_19 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  _T_8679_0_20 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  _T_8679_0_21 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  _T_8679_0_22 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  _T_8679_0_23 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  _T_8679_0_24 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  _T_8679_0_25 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  _T_8679_0_26 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  _T_8679_0_27 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  _T_8679_0_28 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  _T_8679_0_29 = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  _T_8679_0_30 = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  _T_8679_0_31 = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  _T_8898_0 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  _T_8908 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  _T_8911 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  _T_8914 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      if (_T_431) begin
        if (_T_433) begin
          if (_T_435) begin
            _T_239 <= 1'h0;
          end else begin
            _T_239 <= _T_439;
          end
        end
      end
    end
    if (reset) begin
      _T_242 <= 1'h0;
    end else begin
      if (_T_4142) begin
        if (_T_4144) begin
          _T_242 <= 1'h0;
        end else begin
          _T_242 <= _T_4148;
        end
      end
    end
    if (reset) begin
      _T_245 <= 1'h1;
    end else begin
      if (_T_4209) begin
        if (_T_4211) begin
          if (_T_245) begin
            _T_245 <= 1'h1;
          end else begin
            _T_245 <= _T_4217;
          end
        end
      end
    end
    if (reset) begin
      _T_248 <= 1'h1;
    end else begin
      if (_T_7920) begin
        if (_T_248) begin
          _T_248 <= 1'h1;
        end else begin
          _T_248 <= _T_7926;
        end
      end
    end
    if (reset) begin
      _T_251 <= 1'h0;
    end else begin
      if (_T_8522) begin
        if (_T_8525) begin
          if (_T_8527) begin
            _T_251 <= 1'h0;
          end else begin
            _T_251 <= _T_8531;
          end
        end
      end
    end
    if (reset) begin
      _T_254 <= 1'h1;
    end else begin
      if (_T_9121) begin
        if (_T_9124) begin
          if (_T_254) begin
            _T_254 <= 1'h1;
          end else begin
            _T_254 <= _T_9130;
          end
        end
      end
    end
    _T_256 <= cores_0_inputMemAddr;
    _T_258 <= cores_0_inputMemBlockReady;
    _T_260 <= cores_0_inputAddrsIgnore;
    _T_262 <= cores_0_inputBlocksFinished;
    _T_288 <= cores_1_inputMemAddr;
    _T_290 <= cores_1_inputMemBlockReady;
    _T_292 <= cores_1_inputAddrsIgnore;
    _T_294 <= cores_1_inputBlocksFinished;
    _T_320 <= cores_0_outputMemAddr;
    _T_322 <= cores_0_outputMemAddrValid;
    _T_324 <= cores_0_outputMemBlockValid;
    _T_326 <= cores_0_outputMemBlock;
    _T_328 <= cores_0_outputMemIdx;
    _T_330 <= cores_0_outputFinished;
    _T_368 <= cores_1_outputMemAddr;
    _T_370 <= cores_1_outputMemAddrValid;
    _T_372 <= cores_1_outputMemBlockValid;
    _T_374 <= cores_1_outputMemBlock;
    _T_376 <= cores_1_outputMemIdx;
    _T_378 <= cores_1_outputFinished;
    if (reset) begin
      _T_417 <= 1'h0;
    end else begin
      if (_T_431) begin
        if (_T_433) begin
          _T_417 <= 1'h0;
        end else begin
          if (_T_419) begin
            _T_417 <= _T_422;
          end
        end
      end else begin
        if (_T_419) begin
          _T_417 <= _T_422;
        end
      end
    end
    if (reset) begin
      _T_425 <= 1'h0;
    end else begin
      if (_T_431) begin
        if (_T_433) begin
          _T_425 <= 1'h0;
        end else begin
          _T_425 <= _T_445;
        end
      end
    end
    if (reset) begin
      _T_457 <= 1'h0;
    end else begin
      if (_T_4142) begin
        _T_457 <= 1'h0;
      end else begin
        if (_T_459) begin
          _T_457 <= _T_462;
        end
      end
    end
    if (_T_798) begin
      _T_536_0_0 <= _T_902;
    end
    if (_T_798) begin
      _T_536_0_1 <= _T_1006;
    end
    if (_T_798) begin
      _T_536_0_2 <= _T_1110;
    end
    if (_T_798) begin
      _T_536_0_3 <= _T_1214;
    end
    if (_T_798) begin
      _T_536_0_4 <= _T_1318;
    end
    if (_T_798) begin
      _T_536_0_5 <= _T_1422;
    end
    if (_T_798) begin
      _T_536_0_6 <= _T_1526;
    end
    if (_T_798) begin
      _T_536_0_7 <= _T_1630;
    end
    if (_T_798) begin
      _T_536_0_8 <= _T_1734;
    end
    if (_T_798) begin
      _T_536_0_9 <= _T_1838;
    end
    if (_T_798) begin
      _T_536_0_10 <= _T_1942;
    end
    if (_T_798) begin
      _T_536_0_11 <= _T_2046;
    end
    if (_T_798) begin
      _T_536_0_12 <= _T_2150;
    end
    if (_T_798) begin
      _T_536_0_13 <= _T_2254;
    end
    if (_T_798) begin
      _T_536_0_14 <= _T_2358;
    end
    if (_T_798) begin
      _T_536_0_15 <= _T_2462;
    end
    if (_T_798) begin
      _T_536_0_16 <= _T_2566;
    end
    if (_T_798) begin
      _T_536_0_17 <= _T_2670;
    end
    if (_T_798) begin
      _T_536_0_18 <= _T_2774;
    end
    if (_T_798) begin
      _T_536_0_19 <= _T_2878;
    end
    if (_T_798) begin
      _T_536_0_20 <= _T_2982;
    end
    if (_T_798) begin
      _T_536_0_21 <= _T_3086;
    end
    if (_T_798) begin
      _T_536_0_22 <= _T_3190;
    end
    if (_T_798) begin
      _T_536_0_23 <= _T_3294;
    end
    if (_T_798) begin
      _T_536_0_24 <= _T_3398;
    end
    if (_T_798) begin
      _T_536_0_25 <= _T_3502;
    end
    if (_T_798) begin
      _T_536_0_26 <= _T_3606;
    end
    if (_T_798) begin
      _T_536_0_27 <= _T_3710;
    end
    if (_T_798) begin
      _T_536_0_28 <= _T_3814;
    end
    if (_T_798) begin
      _T_536_0_29 <= _T_3918;
    end
    if (_T_798) begin
      _T_536_0_30 <= _T_4022;
    end
    if (_T_798) begin
      _T_536_0_31 <= _T_4126;
    end
    if (reset) begin
      _T_755_0 <= 5'h0;
    end else begin
      if (_T_776_0) begin
        if (_T_4158) begin
          _T_755_0 <= 5'h0;
        end else begin
          _T_755_0 <= _T_4163;
        end
      end
    end
    if (reset) begin
      _T_776_0 <= 1'h0;
    end else begin
      if (_T_776_0) begin
        if (_T_4158) begin
          _T_776_0 <= 1'h0;
        end else begin
          if (_T_798) begin
            _T_776_0 <= _T_4134;
          end
        end
      end else begin
        if (_T_798) begin
          _T_776_0 <= _T_4134;
        end
      end
    end
    if (reset) begin
      _T_786 <= 1'h0;
    end else begin
      if (_T_4142) begin
        _T_786 <= 1'h0;
      end else begin
        if (_T_798) begin
          _T_786 <= _T_4137;
        end
      end
    end
    if (reset) begin
      _T_4195 <= 1'h0;
    end else begin
      if (_T_4209) begin
        if (_T_4211) begin
          _T_4195 <= 1'h0;
        end else begin
          if (_T_4197) begin
            _T_4195 <= _T_4200;
          end
        end
      end else begin
        if (_T_4197) begin
          _T_4195 <= _T_4200;
        end
      end
    end
    if (reset) begin
      _T_4203 <= 1'h0;
    end else begin
      if (_T_4209) begin
        if (_T_4211) begin
          _T_4203 <= 1'h0;
        end else begin
          _T_4203 <= _T_4223;
        end
      end
    end
    if (reset) begin
      _T_4235 <= 1'h0;
    end else begin
      if (_T_7920) begin
        _T_4235 <= 1'h0;
      end else begin
        if (_T_4237) begin
          _T_4235 <= _T_4240;
        end
      end
    end
    if (_T_4576) begin
      _T_4314_0_0 <= _T_4680;
    end
    if (_T_4576) begin
      _T_4314_0_1 <= _T_4784;
    end
    if (_T_4576) begin
      _T_4314_0_2 <= _T_4888;
    end
    if (_T_4576) begin
      _T_4314_0_3 <= _T_4992;
    end
    if (_T_4576) begin
      _T_4314_0_4 <= _T_5096;
    end
    if (_T_4576) begin
      _T_4314_0_5 <= _T_5200;
    end
    if (_T_4576) begin
      _T_4314_0_6 <= _T_5304;
    end
    if (_T_4576) begin
      _T_4314_0_7 <= _T_5408;
    end
    if (_T_4576) begin
      _T_4314_0_8 <= _T_5512;
    end
    if (_T_4576) begin
      _T_4314_0_9 <= _T_5616;
    end
    if (_T_4576) begin
      _T_4314_0_10 <= _T_5720;
    end
    if (_T_4576) begin
      _T_4314_0_11 <= _T_5824;
    end
    if (_T_4576) begin
      _T_4314_0_12 <= _T_5928;
    end
    if (_T_4576) begin
      _T_4314_0_13 <= _T_6032;
    end
    if (_T_4576) begin
      _T_4314_0_14 <= _T_6136;
    end
    if (_T_4576) begin
      _T_4314_0_15 <= _T_6240;
    end
    if (_T_4576) begin
      _T_4314_0_16 <= _T_6344;
    end
    if (_T_4576) begin
      _T_4314_0_17 <= _T_6448;
    end
    if (_T_4576) begin
      _T_4314_0_18 <= _T_6552;
    end
    if (_T_4576) begin
      _T_4314_0_19 <= _T_6656;
    end
    if (_T_4576) begin
      _T_4314_0_20 <= _T_6760;
    end
    if (_T_4576) begin
      _T_4314_0_21 <= _T_6864;
    end
    if (_T_4576) begin
      _T_4314_0_22 <= _T_6968;
    end
    if (_T_4576) begin
      _T_4314_0_23 <= _T_7072;
    end
    if (_T_4576) begin
      _T_4314_0_24 <= _T_7176;
    end
    if (_T_4576) begin
      _T_4314_0_25 <= _T_7280;
    end
    if (_T_4576) begin
      _T_4314_0_26 <= _T_7384;
    end
    if (_T_4576) begin
      _T_4314_0_27 <= _T_7488;
    end
    if (_T_4576) begin
      _T_4314_0_28 <= _T_7592;
    end
    if (_T_4576) begin
      _T_4314_0_29 <= _T_7696;
    end
    if (_T_4576) begin
      _T_4314_0_30 <= _T_7800;
    end
    if (_T_4576) begin
      _T_4314_0_31 <= _T_7904;
    end
    if (reset) begin
      _T_4533_0 <= 5'h0;
    end else begin
      if (_T_4554_0) begin
        if (_T_7936) begin
          _T_4533_0 <= 5'h0;
        end else begin
          _T_4533_0 <= _T_7941;
        end
      end
    end
    if (reset) begin
      _T_4554_0 <= 1'h0;
    end else begin
      if (_T_4554_0) begin
        if (_T_7936) begin
          _T_4554_0 <= 1'h0;
        end else begin
          if (_T_4576) begin
            _T_4554_0 <= _T_7912;
          end
        end
      end else begin
        if (_T_4576) begin
          _T_4554_0 <= _T_7912;
        end
      end
    end
    if (reset) begin
      _T_4564 <= 1'h0;
    end else begin
      if (_T_7920) begin
        _T_4564 <= 1'h0;
      end else begin
        if (_T_4576) begin
          _T_4564 <= _T_7915;
        end
      end
    end
    if (reset) begin
      _T_7973 <= 1'h0;
    end else begin
      if (_T_8522) begin
        if (_T_8525) begin
          _T_7973 <= 1'h0;
        end else begin
          if (_T_7975) begin
            _T_7973 <= _T_7978;
          end
        end
      end else begin
        if (_T_7975) begin
          _T_7973 <= _T_7978;
        end
      end
    end
    if (reset) begin
      _T_7992_0 <= 1'h0;
    end else begin
      if (_T_8522) begin
        if (_T_8525) begin
          _T_7992_0 <= 1'h0;
        end else begin
          if (_T_8342) begin
            _T_7992_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_8342) begin
          _T_7992_0 <= 1'h1;
        end
      end
    end
    if (_T_8342) begin
      _T_8003_0 <= _T_333_0;
    end
    if (_T_345_0) begin
      if (5'h0 == _T_357_0) begin
        _T_8080_0_0 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h1 == _T_357_0) begin
        _T_8080_0_1 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h2 == _T_357_0) begin
        _T_8080_0_2 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h3 == _T_357_0) begin
        _T_8080_0_3 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h4 == _T_357_0) begin
        _T_8080_0_4 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h5 == _T_357_0) begin
        _T_8080_0_5 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h6 == _T_357_0) begin
        _T_8080_0_6 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h7 == _T_357_0) begin
        _T_8080_0_7 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h8 == _T_357_0) begin
        _T_8080_0_8 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h9 == _T_357_0) begin
        _T_8080_0_9 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'ha == _T_357_0) begin
        _T_8080_0_10 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'hb == _T_357_0) begin
        _T_8080_0_11 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'hc == _T_357_0) begin
        _T_8080_0_12 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'hd == _T_357_0) begin
        _T_8080_0_13 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'he == _T_357_0) begin
        _T_8080_0_14 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'hf == _T_357_0) begin
        _T_8080_0_15 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h10 == _T_357_0) begin
        _T_8080_0_16 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h11 == _T_357_0) begin
        _T_8080_0_17 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h12 == _T_357_0) begin
        _T_8080_0_18 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h13 == _T_357_0) begin
        _T_8080_0_19 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h14 == _T_357_0) begin
        _T_8080_0_20 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h15 == _T_357_0) begin
        _T_8080_0_21 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h16 == _T_357_0) begin
        _T_8080_0_22 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h17 == _T_357_0) begin
        _T_8080_0_23 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h18 == _T_357_0) begin
        _T_8080_0_24 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h19 == _T_357_0) begin
        _T_8080_0_25 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h1a == _T_357_0) begin
        _T_8080_0_26 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h1b == _T_357_0) begin
        _T_8080_0_27 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h1c == _T_357_0) begin
        _T_8080_0_28 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h1d == _T_357_0) begin
        _T_8080_0_29 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h1e == _T_357_0) begin
        _T_8080_0_30 <= _GEN_2;
      end
    end
    if (_T_345_0) begin
      if (5'h1f == _T_357_0) begin
        _T_8080_0_31 <= _GEN_2;
      end
    end
    if (reset) begin
      _T_8299_0 <= 1'h0;
    end else begin
      if (_T_8522) begin
        if (_T_8525) begin
          _T_8299_0 <= 1'h0;
        end else begin
          if (_T_8327) begin
            _T_8299_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_8327) begin
          _T_8299_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_8309 <= 1'h0;
    end else begin
      if (_T_8522) begin
        if (_T_8525) begin
          _T_8309 <= 1'h0;
        end else begin
          _T_8309 <= _T_8540;
        end
      end
    end
    if (reset) begin
      _T_8312 <= 1'h0;
    end else begin
      if (_T_8522) begin
        _T_8312 <= 1'h0;
      end else begin
        if (_T_8511) begin
          _T_8312 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_8315 <= 1'h0;
    end else begin
      if (_T_8522) begin
        if (_T_8525) begin
          _T_8315 <= 1'h0;
        end else begin
          if (_T_8320) begin
            _T_8315 <= 1'h1;
          end
        end
      end else begin
        if (_T_8320) begin
          _T_8315 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_8572 <= 1'h0;
    end else begin
      if (_T_9121) begin
        if (_T_9124) begin
          _T_8572 <= 1'h0;
        end else begin
          if (_T_8574) begin
            _T_8572 <= _T_8577;
          end
        end
      end else begin
        if (_T_8574) begin
          _T_8572 <= _T_8577;
        end
      end
    end
    if (reset) begin
      _T_8591_0 <= 1'h0;
    end else begin
      if (_T_9121) begin
        if (_T_9124) begin
          _T_8591_0 <= 1'h0;
        end else begin
          if (_T_8941) begin
            _T_8591_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_8941) begin
          _T_8591_0 <= 1'h1;
        end
      end
    end
    if (_T_8941) begin
      _T_8602_0 <= _T_381_0;
    end
    if (_T_393_0) begin
      if (5'h0 == _T_405_0) begin
        _T_8679_0_0 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h1 == _T_405_0) begin
        _T_8679_0_1 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h2 == _T_405_0) begin
        _T_8679_0_2 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h3 == _T_405_0) begin
        _T_8679_0_3 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h4 == _T_405_0) begin
        _T_8679_0_4 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h5 == _T_405_0) begin
        _T_8679_0_5 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h6 == _T_405_0) begin
        _T_8679_0_6 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h7 == _T_405_0) begin
        _T_8679_0_7 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h8 == _T_405_0) begin
        _T_8679_0_8 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h9 == _T_405_0) begin
        _T_8679_0_9 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'ha == _T_405_0) begin
        _T_8679_0_10 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'hb == _T_405_0) begin
        _T_8679_0_11 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'hc == _T_405_0) begin
        _T_8679_0_12 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'hd == _T_405_0) begin
        _T_8679_0_13 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'he == _T_405_0) begin
        _T_8679_0_14 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'hf == _T_405_0) begin
        _T_8679_0_15 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h10 == _T_405_0) begin
        _T_8679_0_16 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h11 == _T_405_0) begin
        _T_8679_0_17 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h12 == _T_405_0) begin
        _T_8679_0_18 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h13 == _T_405_0) begin
        _T_8679_0_19 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h14 == _T_405_0) begin
        _T_8679_0_20 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h15 == _T_405_0) begin
        _T_8679_0_21 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h16 == _T_405_0) begin
        _T_8679_0_22 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h17 == _T_405_0) begin
        _T_8679_0_23 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h18 == _T_405_0) begin
        _T_8679_0_24 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h19 == _T_405_0) begin
        _T_8679_0_25 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h1a == _T_405_0) begin
        _T_8679_0_26 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h1b == _T_405_0) begin
        _T_8679_0_27 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h1c == _T_405_0) begin
        _T_8679_0_28 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h1d == _T_405_0) begin
        _T_8679_0_29 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h1e == _T_405_0) begin
        _T_8679_0_30 <= _GEN_3;
      end
    end
    if (_T_393_0) begin
      if (5'h1f == _T_405_0) begin
        _T_8679_0_31 <= _GEN_3;
      end
    end
    if (reset) begin
      _T_8898_0 <= 1'h0;
    end else begin
      if (_T_9121) begin
        if (_T_9124) begin
          _T_8898_0 <= 1'h0;
        end else begin
          if (_T_8926) begin
            _T_8898_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_8926) begin
          _T_8898_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_8908 <= 1'h0;
    end else begin
      if (_T_9121) begin
        if (_T_9124) begin
          _T_8908 <= 1'h0;
        end else begin
          _T_8908 <= _T_9139;
        end
      end
    end
    if (reset) begin
      _T_8911 <= 1'h0;
    end else begin
      if (_T_9121) begin
        _T_8911 <= 1'h0;
      end else begin
        if (_T_9110) begin
          _T_8911 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_8914 <= 1'h0;
    end else begin
      if (_T_9121) begin
        if (_T_9124) begin
          _T_8914 <= 1'h0;
        end else begin
          if (_T_8919) begin
            _T_8914 <= 1'h1;
          end
        end
      end else begin
        if (_T_8919) begin
          _T_8914 <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_794 & _T_4156) begin
          $fwrite(32'h80000002,"inputBuffer: 0x%h for core %d, channel 0\n",io_inputMemBlocks_0,_T_4153);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4572 & _T_4156) begin
          $fwrite(32'h80000002,"inputBuffer: 0x%h for core %d, channel 1\n",io_inputMemBlocks_1,_T_7931);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8565 & _T_4156) begin
          $fwrite(32'h80000002,"outputBuffer: 0x%h for core %d, channel 0\n",io_outputMemBlocks_0,_T_8566);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9164 & _T_4156) begin
          $fwrite(32'h80000002,"outputBuffer: 0x%h for core %d, channel 1\n",io_outputMemBlocks_1,_T_9165);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
