`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module StreamingMemoryController(
  input          clock,
  input          reset,
  output [63:0]  io_axi_inputMemAddrs_0,
  output [63:0]  io_axi_inputMemAddrs_1,
  output [63:0]  io_axi_inputMemAddrs_2,
  output [63:0]  io_axi_inputMemAddrs_3,
  output         io_axi_inputMemAddrValids_0,
  output         io_axi_inputMemAddrValids_1,
  output         io_axi_inputMemAddrValids_2,
  output         io_axi_inputMemAddrValids_3,
  output [7:0]   io_axi_inputMemAddrLens_0,
  output [7:0]   io_axi_inputMemAddrLens_1,
  output [7:0]   io_axi_inputMemAddrLens_2,
  output [7:0]   io_axi_inputMemAddrLens_3,
  input          io_axi_inputMemAddrReadys_0,
  input          io_axi_inputMemAddrReadys_1,
  input          io_axi_inputMemAddrReadys_2,
  input          io_axi_inputMemAddrReadys_3,
  input  [511:0] io_axi_inputMemBlocks_0,
  input  [511:0] io_axi_inputMemBlocks_1,
  input  [511:0] io_axi_inputMemBlocks_2,
  input  [511:0] io_axi_inputMemBlocks_3,
  input          io_axi_inputMemBlockValids_0,
  input          io_axi_inputMemBlockValids_1,
  input          io_axi_inputMemBlockValids_2,
  input          io_axi_inputMemBlockValids_3,
  output         io_axi_inputMemBlockReadys_0,
  output         io_axi_inputMemBlockReadys_1,
  output         io_axi_inputMemBlockReadys_2,
  output         io_axi_inputMemBlockReadys_3,
  output [63:0]  io_axi_outputMemAddrs_0,
  output [63:0]  io_axi_outputMemAddrs_1,
  output [63:0]  io_axi_outputMemAddrs_2,
  output [63:0]  io_axi_outputMemAddrs_3,
  output         io_axi_outputMemAddrValids_0,
  output         io_axi_outputMemAddrValids_1,
  output         io_axi_outputMemAddrValids_2,
  output         io_axi_outputMemAddrValids_3,
  output [7:0]   io_axi_outputMemAddrLens_0,
  output [7:0]   io_axi_outputMemAddrLens_1,
  output [7:0]   io_axi_outputMemAddrLens_2,
  output [7:0]   io_axi_outputMemAddrLens_3,
  output [15:0]  io_axi_outputMemAddrIds_0,
  output [15:0]  io_axi_outputMemAddrIds_1,
  output [15:0]  io_axi_outputMemAddrIds_2,
  output [15:0]  io_axi_outputMemAddrIds_3,
  input          io_axi_outputMemAddrReadys_0,
  input          io_axi_outputMemAddrReadys_1,
  input          io_axi_outputMemAddrReadys_2,
  input          io_axi_outputMemAddrReadys_3,
  output [511:0] io_axi_outputMemBlocks_0,
  output [511:0] io_axi_outputMemBlocks_1,
  output [511:0] io_axi_outputMemBlocks_2,
  output [511:0] io_axi_outputMemBlocks_3,
  output         io_axi_outputMemBlockValids_0,
  output         io_axi_outputMemBlockValids_1,
  output         io_axi_outputMemBlockValids_2,
  output         io_axi_outputMemBlockValids_3,
  output         io_axi_outputMemBlockLasts_0,
  output         io_axi_outputMemBlockLasts_1,
  output         io_axi_outputMemBlockLasts_2,
  output         io_axi_outputMemBlockLasts_3,
  input          io_axi_outputMemBlockReadys_0,
  input          io_axi_outputMemBlockReadys_1,
  input          io_axi_outputMemBlockReadys_2,
  input          io_axi_outputMemBlockReadys_3,
  output         io_axi_finished,
  output [31:0]  io_streamingCores_0_metadataPtr,
  input  [31:0]  io_streamingCores_0_inputMemAddr,
  input          io_streamingCores_0_inputMemAddrValid,
  input          io_streamingCores_0_inputMemAddrsFinished,
  output [31:0]  io_streamingCores_0_inputMemBlock,
  output [4:0]   io_streamingCores_0_inputMemIdx,
  output         io_streamingCores_0_inputMemBlockValid,
  input  [31:0]  io_streamingCores_0_outputMemAddr,
  input          io_streamingCores_0_outputMemAddrValid,
  output         io_streamingCores_0_outputMemAddrReady,
  input  [31:0]  io_streamingCores_0_outputMemBlock,
  input  [4:0]   io_streamingCores_0_outputMemIdx,
  input          io_streamingCores_0_outputMemBlockValid,
  input          io_streamingCores_0_outputFinished,
  output [31:0]  io_streamingCores_1_metadataPtr,
  input  [31:0]  io_streamingCores_1_inputMemAddr,
  input          io_streamingCores_1_inputMemAddrValid,
  input          io_streamingCores_1_inputMemAddrsFinished,
  output [31:0]  io_streamingCores_1_inputMemBlock,
  output [4:0]   io_streamingCores_1_inputMemIdx,
  output         io_streamingCores_1_inputMemBlockValid,
  input  [31:0]  io_streamingCores_1_outputMemAddr,
  input          io_streamingCores_1_outputMemAddrValid,
  output         io_streamingCores_1_outputMemAddrReady,
  input  [31:0]  io_streamingCores_1_outputMemBlock,
  input  [4:0]   io_streamingCores_1_outputMemIdx,
  input          io_streamingCores_1_outputMemBlockValid,
  input          io_streamingCores_1_outputFinished,
  output [31:0]  io_streamingCores_2_metadataPtr,
  input  [31:0]  io_streamingCores_2_inputMemAddr,
  input          io_streamingCores_2_inputMemAddrValid,
  input          io_streamingCores_2_inputMemAddrsFinished,
  output [31:0]  io_streamingCores_2_inputMemBlock,
  output [4:0]   io_streamingCores_2_inputMemIdx,
  output         io_streamingCores_2_inputMemBlockValid,
  input  [31:0]  io_streamingCores_2_outputMemAddr,
  input          io_streamingCores_2_outputMemAddrValid,
  output         io_streamingCores_2_outputMemAddrReady,
  input  [31:0]  io_streamingCores_2_outputMemBlock,
  input  [4:0]   io_streamingCores_2_outputMemIdx,
  input          io_streamingCores_2_outputMemBlockValid,
  input          io_streamingCores_2_outputFinished,
  output [31:0]  io_streamingCores_3_metadataPtr,
  input  [31:0]  io_streamingCores_3_inputMemAddr,
  input          io_streamingCores_3_inputMemAddrValid,
  input          io_streamingCores_3_inputMemAddrsFinished,
  output [31:0]  io_streamingCores_3_inputMemBlock,
  output [4:0]   io_streamingCores_3_inputMemIdx,
  output         io_streamingCores_3_inputMemBlockValid,
  input  [31:0]  io_streamingCores_3_outputMemAddr,
  input          io_streamingCores_3_outputMemAddrValid,
  output         io_streamingCores_3_outputMemAddrReady,
  input  [31:0]  io_streamingCores_3_outputMemBlock,
  input  [4:0]   io_streamingCores_3_outputMemIdx,
  input          io_streamingCores_3_outputMemBlockValid,
  input          io_streamingCores_3_outputFinished
);
  reg  _T_389;
  reg [31:0] _RAND_0;
  reg  _T_395;
  reg [31:0] _RAND_1;
  reg  _T_401;
  reg [31:0] _RAND_2;
  reg  _T_407;
  reg [31:0] _RAND_3;
  reg  _T_410;
  reg [31:0] _RAND_4;
  reg  _T_413;
  reg [31:0] _RAND_5;
  reg  _T_416;
  reg [31:0] _RAND_6;
  reg  _T_419;
  reg [31:0] _RAND_7;
  wire [31:0] _T_422_0;
  wire  _T_428_0;
  wire  _T_434_0;
  wire [31:0] _T_440_0;
  wire  _T_446_0;
  wire  _T_452_0;
  wire [31:0] _T_458_0;
  wire  _T_464_0;
  wire  _T_470_0;
  wire [31:0] _T_476_0;
  wire  _T_482_0;
  wire  _T_488_0;
  wire [31:0] _T_494_0;
  wire  _T_500_0;
  wire  _T_506_0;
  wire [31:0] _T_512_0;
  wire [4:0] _T_518_0;
  wire  _T_524_0;
  wire [31:0] _T_530_0;
  wire  _T_536_0;
  wire  _T_542_0;
  wire [31:0] _T_548_0;
  wire [4:0] _T_554_0;
  wire  _T_560_0;
  wire [31:0] _T_566_0;
  wire  _T_572_0;
  wire  _T_578_0;
  wire [31:0] _T_584_0;
  wire [4:0] _T_590_0;
  wire  _T_596_0;
  wire [31:0] _T_602_0;
  wire  _T_608_0;
  wire  _T_614_0;
  wire [31:0] _T_620_0;
  wire [4:0] _T_626_0;
  wire  _T_632_0;
  reg  _T_638;
  reg [31:0] _RAND_8;
  reg  _T_652_0;
  reg [31:0] _RAND_9;
  reg  _T_673_0;
  reg [31:0] _RAND_10;
  reg [31:0] _T_754_0_0;
  reg [31:0] _RAND_11;
  reg [31:0] _T_754_0_1;
  reg [31:0] _RAND_12;
  reg [31:0] _T_754_0_2;
  reg [31:0] _RAND_13;
  reg [31:0] _T_754_0_3;
  reg [31:0] _RAND_14;
  reg [31:0] _T_754_0_4;
  reg [31:0] _RAND_15;
  reg [31:0] _T_754_0_5;
  reg [31:0] _RAND_16;
  reg [31:0] _T_754_0_6;
  reg [31:0] _RAND_17;
  reg [31:0] _T_754_0_7;
  reg [31:0] _RAND_18;
  reg [31:0] _T_754_0_8;
  reg [31:0] _RAND_19;
  reg [31:0] _T_754_0_9;
  reg [31:0] _RAND_20;
  reg [31:0] _T_754_0_10;
  reg [31:0] _RAND_21;
  reg [31:0] _T_754_0_11;
  reg [31:0] _RAND_22;
  reg [31:0] _T_754_0_12;
  reg [31:0] _RAND_23;
  reg [31:0] _T_754_0_13;
  reg [31:0] _RAND_24;
  reg [31:0] _T_754_0_14;
  reg [31:0] _RAND_25;
  reg [31:0] _T_754_0_15;
  reg [31:0] _RAND_26;
  reg [31:0] _T_754_0_16;
  reg [31:0] _RAND_27;
  reg [31:0] _T_754_0_17;
  reg [31:0] _RAND_28;
  reg [31:0] _T_754_0_18;
  reg [31:0] _RAND_29;
  reg [31:0] _T_754_0_19;
  reg [31:0] _RAND_30;
  reg [31:0] _T_754_0_20;
  reg [31:0] _RAND_31;
  reg [31:0] _T_754_0_21;
  reg [31:0] _RAND_32;
  reg [31:0] _T_754_0_22;
  reg [31:0] _RAND_33;
  reg [31:0] _T_754_0_23;
  reg [31:0] _RAND_34;
  reg [31:0] _T_754_0_24;
  reg [31:0] _RAND_35;
  reg [31:0] _T_754_0_25;
  reg [31:0] _RAND_36;
  reg [31:0] _T_754_0_26;
  reg [31:0] _RAND_37;
  reg [31:0] _T_754_0_27;
  reg [31:0] _RAND_38;
  reg [31:0] _T_754_0_28;
  reg [31:0] _RAND_39;
  reg [31:0] _T_754_0_29;
  reg [31:0] _RAND_40;
  reg [31:0] _T_754_0_30;
  reg [31:0] _RAND_41;
  reg [31:0] _T_754_0_31;
  reg [31:0] _RAND_42;
  reg [4:0] _T_973_0;
  reg [31:0] _RAND_43;
  reg  _T_994_0;
  reg [31:0] _RAND_44;
  reg  _T_1004;
  reg [31:0] _RAND_45;
  reg  _T_1007;
  reg [31:0] _RAND_46;
  reg  _T_1010;
  reg [31:0] _RAND_47;
  wire  _T_1014;
  wire  _T_1016;
  wire [1:0] _T_1018;
  wire  _T_1019;
  wire  _GEN_8;
  wire  _T_1026;
  wire  _T_1032;
  wire  _T_1033;
  wire  _T_1035;
  wire  _T_1040;
  wire  _T_1047;
  wire  _T_1048;
  wire  _GEN_9;
  wire  _T_1060;
  wire [1:0] _T_1071;
  wire  _T_1072;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _T_1074;
  wire [5:0] _T_1080;
  wire [4:0] _T_1081;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire [4:0] _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire  _GEN_24;
  wire [4:0] _GEN_25;
  wire  _T_1082;
  wire [1:0] _T_1087;
  wire  _T_1088;
  wire  _T_1089;
  wire  _T_1091;
  wire [31:0] _T_1195;
  wire [31:0] _GEN_26;
  wire [31:0] _T_1301;
  wire [31:0] _GEN_27;
  wire [31:0] _T_1407;
  wire [31:0] _GEN_28;
  wire [31:0] _T_1513;
  wire [31:0] _GEN_29;
  wire [31:0] _T_1619;
  wire [31:0] _GEN_30;
  wire [31:0] _T_1725;
  wire [31:0] _GEN_31;
  wire [31:0] _T_1831;
  wire [31:0] _GEN_32;
  wire [31:0] _T_1937;
  wire [31:0] _GEN_33;
  wire [31:0] _T_2043;
  wire [31:0] _GEN_34;
  wire [31:0] _T_2149;
  wire [31:0] _GEN_35;
  wire [31:0] _T_2255;
  wire [31:0] _GEN_36;
  wire [31:0] _T_2361;
  wire [31:0] _GEN_37;
  wire [31:0] _T_2467;
  wire [31:0] _GEN_38;
  wire [31:0] _T_2573;
  wire [31:0] _GEN_39;
  wire [31:0] _T_2679;
  wire [31:0] _GEN_40;
  wire [31:0] _T_2785;
  wire [31:0] _GEN_41;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  wire [31:0] _GEN_44;
  wire [31:0] _GEN_45;
  wire [31:0] _GEN_46;
  wire [31:0] _GEN_47;
  wire [31:0] _GEN_48;
  wire [31:0] _GEN_49;
  wire [31:0] _GEN_50;
  wire [31:0] _GEN_51;
  wire [31:0] _GEN_52;
  wire [31:0] _GEN_53;
  wire [31:0] _GEN_54;
  wire [31:0] _GEN_55;
  wire [31:0] _GEN_56;
  wire [31:0] _GEN_57;
  wire  _GEN_58;
  wire [31:0] _GEN_59;
  wire [31:0] _GEN_60;
  wire [31:0] _GEN_61;
  wire [31:0] _GEN_62;
  wire [31:0] _GEN_63;
  wire [31:0] _GEN_64;
  wire [31:0] _GEN_65;
  wire [31:0] _GEN_66;
  wire [31:0] _GEN_67;
  wire [31:0] _GEN_68;
  wire [31:0] _GEN_69;
  wire [31:0] _GEN_70;
  wire [31:0] _GEN_71;
  wire [31:0] _GEN_72;
  wire [31:0] _GEN_73;
  wire [31:0] _GEN_74;
  wire [31:0] _GEN_75;
  wire [31:0] _GEN_76;
  wire [31:0] _GEN_77;
  wire [31:0] _GEN_78;
  wire [31:0] _GEN_79;
  wire [31:0] _GEN_80;
  wire [31:0] _GEN_81;
  wire [31:0] _GEN_82;
  wire [31:0] _GEN_83;
  wire [31:0] _GEN_84;
  wire [31:0] _GEN_85;
  wire [31:0] _GEN_86;
  wire [31:0] _GEN_87;
  wire [31:0] _GEN_88;
  wire [31:0] _GEN_89;
  wire [31:0] _GEN_90;
  wire  _T_4482;
  wire  _T_4485;
  wire  _T_4495;
  wire  _T_4496;
  wire  _T_4502;
  wire  _T_4503;
  wire  _T_4504;
  wire  _GEN_91;
  wire  _GEN_92;
  wire  _T_4516;
  wire  _T_4518;
  wire [1:0] _T_4521;
  wire  _T_4522;
  wire  _T_4523;
  wire [1:0] _T_4526;
  wire  _T_4527;
  wire  _GEN_93;
  wire  _GEN_94;
  wire  _GEN_95;
  wire  _GEN_96;
  wire  _GEN_97;
  wire  _GEN_98;
  wire  _T_4538;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_99;
  wire [31:0] _GEN_100;
  wire [31:0] _GEN_101;
  wire [31:0] _GEN_102;
  wire [31:0] _GEN_103;
  wire [31:0] _GEN_104;
  wire [31:0] _GEN_105;
  wire [31:0] _GEN_106;
  wire [31:0] _GEN_107;
  wire [31:0] _GEN_108;
  wire [31:0] _GEN_109;
  wire [31:0] _GEN_110;
  wire [31:0] _GEN_111;
  wire [31:0] _GEN_112;
  wire [31:0] _GEN_113;
  wire [31:0] _GEN_114;
  wire [31:0] _GEN_115;
  wire [31:0] _GEN_116;
  wire [31:0] _GEN_117;
  wire [31:0] _GEN_118;
  wire [31:0] _GEN_119;
  wire [31:0] _GEN_120;
  wire [31:0] _GEN_121;
  wire [31:0] _GEN_122;
  wire [31:0] _GEN_123;
  wire [31:0] _GEN_124;
  wire [31:0] _GEN_125;
  wire [31:0] _GEN_126;
  wire [31:0] _GEN_127;
  wire [31:0] _GEN_128;
  wire [31:0] _GEN_129;
  wire [1:0] _T_4545;
  wire [1:0] _T_4546;
  wire  _T_4547;
  wire  _T_4548;
  wire  _T_4550;
  wire  _T_4551;
  wire  _T_4553;
  wire  _T_4555;
  reg  _T_4558;
  reg [31:0] _RAND_48;
  reg  _T_4572_0;
  reg [31:0] _RAND_49;
  reg  _T_4593_0;
  reg [31:0] _RAND_50;
  reg [31:0] _T_4674_0_0;
  reg [31:0] _RAND_51;
  reg [31:0] _T_4674_0_1;
  reg [31:0] _RAND_52;
  reg [31:0] _T_4674_0_2;
  reg [31:0] _RAND_53;
  reg [31:0] _T_4674_0_3;
  reg [31:0] _RAND_54;
  reg [31:0] _T_4674_0_4;
  reg [31:0] _RAND_55;
  reg [31:0] _T_4674_0_5;
  reg [31:0] _RAND_56;
  reg [31:0] _T_4674_0_6;
  reg [31:0] _RAND_57;
  reg [31:0] _T_4674_0_7;
  reg [31:0] _RAND_58;
  reg [31:0] _T_4674_0_8;
  reg [31:0] _RAND_59;
  reg [31:0] _T_4674_0_9;
  reg [31:0] _RAND_60;
  reg [31:0] _T_4674_0_10;
  reg [31:0] _RAND_61;
  reg [31:0] _T_4674_0_11;
  reg [31:0] _RAND_62;
  reg [31:0] _T_4674_0_12;
  reg [31:0] _RAND_63;
  reg [31:0] _T_4674_0_13;
  reg [31:0] _RAND_64;
  reg [31:0] _T_4674_0_14;
  reg [31:0] _RAND_65;
  reg [31:0] _T_4674_0_15;
  reg [31:0] _RAND_66;
  reg [31:0] _T_4674_0_16;
  reg [31:0] _RAND_67;
  reg [31:0] _T_4674_0_17;
  reg [31:0] _RAND_68;
  reg [31:0] _T_4674_0_18;
  reg [31:0] _RAND_69;
  reg [31:0] _T_4674_0_19;
  reg [31:0] _RAND_70;
  reg [31:0] _T_4674_0_20;
  reg [31:0] _RAND_71;
  reg [31:0] _T_4674_0_21;
  reg [31:0] _RAND_72;
  reg [31:0] _T_4674_0_22;
  reg [31:0] _RAND_73;
  reg [31:0] _T_4674_0_23;
  reg [31:0] _RAND_74;
  reg [31:0] _T_4674_0_24;
  reg [31:0] _RAND_75;
  reg [31:0] _T_4674_0_25;
  reg [31:0] _RAND_76;
  reg [31:0] _T_4674_0_26;
  reg [31:0] _RAND_77;
  reg [31:0] _T_4674_0_27;
  reg [31:0] _RAND_78;
  reg [31:0] _T_4674_0_28;
  reg [31:0] _RAND_79;
  reg [31:0] _T_4674_0_29;
  reg [31:0] _RAND_80;
  reg [31:0] _T_4674_0_30;
  reg [31:0] _RAND_81;
  reg [31:0] _T_4674_0_31;
  reg [31:0] _RAND_82;
  reg [4:0] _T_4893_0;
  reg [31:0] _RAND_83;
  reg  _T_4914_0;
  reg [31:0] _RAND_84;
  reg  _T_4924;
  reg [31:0] _RAND_85;
  reg  _T_4927;
  reg [31:0] _RAND_86;
  reg  _T_4930;
  reg [31:0] _RAND_87;
  wire  _T_4934;
  wire  _T_4936;
  wire [1:0] _T_4938;
  wire  _T_4939;
  wire  _GEN_130;
  wire  _T_4946;
  wire  _T_4952;
  wire  _T_4953;
  wire  _T_4955;
  wire  _T_4960;
  wire  _T_4967;
  wire  _T_4968;
  wire  _GEN_131;
  wire  _T_4980;
  wire [1:0] _T_4991;
  wire  _T_4992;
  wire  _GEN_133;
  wire  _GEN_134;
  wire  _GEN_135;
  wire  _GEN_136;
  wire  _GEN_138;
  wire  _GEN_139;
  wire  _T_4994;
  wire [5:0] _T_5000;
  wire [4:0] _T_5001;
  wire  _GEN_140;
  wire  _GEN_141;
  wire  _GEN_142;
  wire [4:0] _GEN_143;
  wire  _GEN_144;
  wire  _GEN_145;
  wire  _GEN_146;
  wire [4:0] _GEN_147;
  wire  _T_5002;
  wire [1:0] _T_5007;
  wire  _T_5008;
  wire  _T_5009;
  wire  _T_5011;
  wire [31:0] _T_5115;
  wire [31:0] _GEN_148;
  wire [31:0] _T_5221;
  wire [31:0] _GEN_149;
  wire [31:0] _T_5327;
  wire [31:0] _GEN_150;
  wire [31:0] _T_5433;
  wire [31:0] _GEN_151;
  wire [31:0] _T_5539;
  wire [31:0] _GEN_152;
  wire [31:0] _T_5645;
  wire [31:0] _GEN_153;
  wire [31:0] _T_5751;
  wire [31:0] _GEN_154;
  wire [31:0] _T_5857;
  wire [31:0] _GEN_155;
  wire [31:0] _T_5963;
  wire [31:0] _GEN_156;
  wire [31:0] _T_6069;
  wire [31:0] _GEN_157;
  wire [31:0] _T_6175;
  wire [31:0] _GEN_158;
  wire [31:0] _T_6281;
  wire [31:0] _GEN_159;
  wire [31:0] _T_6387;
  wire [31:0] _GEN_160;
  wire [31:0] _T_6493;
  wire [31:0] _GEN_161;
  wire [31:0] _T_6599;
  wire [31:0] _GEN_162;
  wire [31:0] _T_6705;
  wire [31:0] _GEN_163;
  wire [31:0] _GEN_164;
  wire [31:0] _GEN_165;
  wire [31:0] _GEN_166;
  wire [31:0] _GEN_167;
  wire [31:0] _GEN_168;
  wire [31:0] _GEN_169;
  wire [31:0] _GEN_170;
  wire [31:0] _GEN_171;
  wire [31:0] _GEN_172;
  wire [31:0] _GEN_173;
  wire [31:0] _GEN_174;
  wire [31:0] _GEN_175;
  wire [31:0] _GEN_176;
  wire [31:0] _GEN_177;
  wire [31:0] _GEN_178;
  wire [31:0] _GEN_179;
  wire  _GEN_180;
  wire [31:0] _GEN_181;
  wire [31:0] _GEN_182;
  wire [31:0] _GEN_183;
  wire [31:0] _GEN_184;
  wire [31:0] _GEN_185;
  wire [31:0] _GEN_186;
  wire [31:0] _GEN_187;
  wire [31:0] _GEN_188;
  wire [31:0] _GEN_189;
  wire [31:0] _GEN_190;
  wire [31:0] _GEN_191;
  wire [31:0] _GEN_192;
  wire [31:0] _GEN_193;
  wire [31:0] _GEN_194;
  wire [31:0] _GEN_195;
  wire [31:0] _GEN_196;
  wire [31:0] _GEN_197;
  wire [31:0] _GEN_198;
  wire [31:0] _GEN_199;
  wire [31:0] _GEN_200;
  wire [31:0] _GEN_201;
  wire [31:0] _GEN_202;
  wire [31:0] _GEN_203;
  wire [31:0] _GEN_204;
  wire [31:0] _GEN_205;
  wire [31:0] _GEN_206;
  wire [31:0] _GEN_207;
  wire [31:0] _GEN_208;
  wire [31:0] _GEN_209;
  wire [31:0] _GEN_210;
  wire [31:0] _GEN_211;
  wire [31:0] _GEN_212;
  wire  _T_8402;
  wire  _T_8405;
  wire  _T_8415;
  wire  _T_8416;
  wire  _T_8422;
  wire  _T_8423;
  wire  _T_8424;
  wire  _GEN_213;
  wire  _GEN_214;
  wire  _T_8436;
  wire  _T_8438;
  wire [1:0] _T_8441;
  wire  _T_8442;
  wire  _T_8443;
  wire [1:0] _T_8446;
  wire  _T_8447;
  wire  _GEN_215;
  wire  _GEN_216;
  wire  _GEN_217;
  wire  _GEN_218;
  wire  _GEN_219;
  wire  _GEN_220;
  wire  _T_8458;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_221;
  wire [31:0] _GEN_222;
  wire [31:0] _GEN_223;
  wire [31:0] _GEN_224;
  wire [31:0] _GEN_225;
  wire [31:0] _GEN_226;
  wire [31:0] _GEN_227;
  wire [31:0] _GEN_228;
  wire [31:0] _GEN_229;
  wire [31:0] _GEN_230;
  wire [31:0] _GEN_231;
  wire [31:0] _GEN_232;
  wire [31:0] _GEN_233;
  wire [31:0] _GEN_234;
  wire [31:0] _GEN_235;
  wire [31:0] _GEN_236;
  wire [31:0] _GEN_237;
  wire [31:0] _GEN_238;
  wire [31:0] _GEN_239;
  wire [31:0] _GEN_240;
  wire [31:0] _GEN_241;
  wire [31:0] _GEN_242;
  wire [31:0] _GEN_243;
  wire [31:0] _GEN_244;
  wire [31:0] _GEN_245;
  wire [31:0] _GEN_246;
  wire [31:0] _GEN_247;
  wire [31:0] _GEN_248;
  wire [31:0] _GEN_249;
  wire [31:0] _GEN_250;
  wire [31:0] _GEN_251;
  wire [1:0] _T_8465;
  wire [1:0] _T_8466;
  wire  _T_8467;
  wire  _T_8468;
  wire  _T_8470;
  wire  _T_8471;
  wire  _T_8473;
  wire  _T_8475;
  reg  _T_8478;
  reg [31:0] _RAND_88;
  reg  _T_8492_0;
  reg [31:0] _RAND_89;
  reg  _T_8513_0;
  reg [31:0] _RAND_90;
  reg [31:0] _T_8594_0_0;
  reg [31:0] _RAND_91;
  reg [31:0] _T_8594_0_1;
  reg [31:0] _RAND_92;
  reg [31:0] _T_8594_0_2;
  reg [31:0] _RAND_93;
  reg [31:0] _T_8594_0_3;
  reg [31:0] _RAND_94;
  reg [31:0] _T_8594_0_4;
  reg [31:0] _RAND_95;
  reg [31:0] _T_8594_0_5;
  reg [31:0] _RAND_96;
  reg [31:0] _T_8594_0_6;
  reg [31:0] _RAND_97;
  reg [31:0] _T_8594_0_7;
  reg [31:0] _RAND_98;
  reg [31:0] _T_8594_0_8;
  reg [31:0] _RAND_99;
  reg [31:0] _T_8594_0_9;
  reg [31:0] _RAND_100;
  reg [31:0] _T_8594_0_10;
  reg [31:0] _RAND_101;
  reg [31:0] _T_8594_0_11;
  reg [31:0] _RAND_102;
  reg [31:0] _T_8594_0_12;
  reg [31:0] _RAND_103;
  reg [31:0] _T_8594_0_13;
  reg [31:0] _RAND_104;
  reg [31:0] _T_8594_0_14;
  reg [31:0] _RAND_105;
  reg [31:0] _T_8594_0_15;
  reg [31:0] _RAND_106;
  reg [31:0] _T_8594_0_16;
  reg [31:0] _RAND_107;
  reg [31:0] _T_8594_0_17;
  reg [31:0] _RAND_108;
  reg [31:0] _T_8594_0_18;
  reg [31:0] _RAND_109;
  reg [31:0] _T_8594_0_19;
  reg [31:0] _RAND_110;
  reg [31:0] _T_8594_0_20;
  reg [31:0] _RAND_111;
  reg [31:0] _T_8594_0_21;
  reg [31:0] _RAND_112;
  reg [31:0] _T_8594_0_22;
  reg [31:0] _RAND_113;
  reg [31:0] _T_8594_0_23;
  reg [31:0] _RAND_114;
  reg [31:0] _T_8594_0_24;
  reg [31:0] _RAND_115;
  reg [31:0] _T_8594_0_25;
  reg [31:0] _RAND_116;
  reg [31:0] _T_8594_0_26;
  reg [31:0] _RAND_117;
  reg [31:0] _T_8594_0_27;
  reg [31:0] _RAND_118;
  reg [31:0] _T_8594_0_28;
  reg [31:0] _RAND_119;
  reg [31:0] _T_8594_0_29;
  reg [31:0] _RAND_120;
  reg [31:0] _T_8594_0_30;
  reg [31:0] _RAND_121;
  reg [31:0] _T_8594_0_31;
  reg [31:0] _RAND_122;
  reg [4:0] _T_8813_0;
  reg [31:0] _RAND_123;
  reg  _T_8834_0;
  reg [31:0] _RAND_124;
  reg  _T_8844;
  reg [31:0] _RAND_125;
  reg  _T_8847;
  reg [31:0] _RAND_126;
  reg  _T_8850;
  reg [31:0] _RAND_127;
  wire  _T_8854;
  wire  _T_8856;
  wire [1:0] _T_8858;
  wire  _T_8859;
  wire  _GEN_252;
  wire  _T_8866;
  wire  _T_8872;
  wire  _T_8873;
  wire  _T_8875;
  wire  _T_8880;
  wire  _T_8887;
  wire  _T_8888;
  wire  _GEN_253;
  wire  _T_8900;
  wire [1:0] _T_8911;
  wire  _T_8912;
  wire  _GEN_255;
  wire  _GEN_256;
  wire  _GEN_257;
  wire  _GEN_258;
  wire  _GEN_260;
  wire  _GEN_261;
  wire  _T_8914;
  wire [5:0] _T_8920;
  wire [4:0] _T_8921;
  wire  _GEN_262;
  wire  _GEN_263;
  wire  _GEN_264;
  wire [4:0] _GEN_265;
  wire  _GEN_266;
  wire  _GEN_267;
  wire  _GEN_268;
  wire [4:0] _GEN_269;
  wire  _T_8922;
  wire [1:0] _T_8927;
  wire  _T_8928;
  wire  _T_8929;
  wire  _T_8931;
  wire [31:0] _T_9035;
  wire [31:0] _GEN_270;
  wire [31:0] _T_9141;
  wire [31:0] _GEN_271;
  wire [31:0] _T_9247;
  wire [31:0] _GEN_272;
  wire [31:0] _T_9353;
  wire [31:0] _GEN_273;
  wire [31:0] _T_9459;
  wire [31:0] _GEN_274;
  wire [31:0] _T_9565;
  wire [31:0] _GEN_275;
  wire [31:0] _T_9671;
  wire [31:0] _GEN_276;
  wire [31:0] _T_9777;
  wire [31:0] _GEN_277;
  wire [31:0] _T_9883;
  wire [31:0] _GEN_278;
  wire [31:0] _T_9989;
  wire [31:0] _GEN_279;
  wire [31:0] _T_10095;
  wire [31:0] _GEN_280;
  wire [31:0] _T_10201;
  wire [31:0] _GEN_281;
  wire [31:0] _T_10307;
  wire [31:0] _GEN_282;
  wire [31:0] _T_10413;
  wire [31:0] _GEN_283;
  wire [31:0] _T_10519;
  wire [31:0] _GEN_284;
  wire [31:0] _T_10625;
  wire [31:0] _GEN_285;
  wire [31:0] _GEN_286;
  wire [31:0] _GEN_287;
  wire [31:0] _GEN_288;
  wire [31:0] _GEN_289;
  wire [31:0] _GEN_290;
  wire [31:0] _GEN_291;
  wire [31:0] _GEN_292;
  wire [31:0] _GEN_293;
  wire [31:0] _GEN_294;
  wire [31:0] _GEN_295;
  wire [31:0] _GEN_296;
  wire [31:0] _GEN_297;
  wire [31:0] _GEN_298;
  wire [31:0] _GEN_299;
  wire [31:0] _GEN_300;
  wire [31:0] _GEN_301;
  wire  _GEN_302;
  wire [31:0] _GEN_303;
  wire [31:0] _GEN_304;
  wire [31:0] _GEN_305;
  wire [31:0] _GEN_306;
  wire [31:0] _GEN_307;
  wire [31:0] _GEN_308;
  wire [31:0] _GEN_309;
  wire [31:0] _GEN_310;
  wire [31:0] _GEN_311;
  wire [31:0] _GEN_312;
  wire [31:0] _GEN_313;
  wire [31:0] _GEN_314;
  wire [31:0] _GEN_315;
  wire [31:0] _GEN_316;
  wire [31:0] _GEN_317;
  wire [31:0] _GEN_318;
  wire [31:0] _GEN_319;
  wire [31:0] _GEN_320;
  wire [31:0] _GEN_321;
  wire [31:0] _GEN_322;
  wire [31:0] _GEN_323;
  wire [31:0] _GEN_324;
  wire [31:0] _GEN_325;
  wire [31:0] _GEN_326;
  wire [31:0] _GEN_327;
  wire [31:0] _GEN_328;
  wire [31:0] _GEN_329;
  wire [31:0] _GEN_330;
  wire [31:0] _GEN_331;
  wire [31:0] _GEN_332;
  wire [31:0] _GEN_333;
  wire [31:0] _GEN_334;
  wire  _T_12322;
  wire  _T_12325;
  wire  _T_12335;
  wire  _T_12336;
  wire  _T_12342;
  wire  _T_12343;
  wire  _T_12344;
  wire  _GEN_335;
  wire  _GEN_336;
  wire  _T_12356;
  wire  _T_12358;
  wire [1:0] _T_12361;
  wire  _T_12362;
  wire  _T_12363;
  wire [1:0] _T_12366;
  wire  _T_12367;
  wire  _GEN_337;
  wire  _GEN_338;
  wire  _GEN_339;
  wire  _GEN_340;
  wire  _GEN_341;
  wire  _GEN_342;
  wire  _T_12378;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_343;
  wire [31:0] _GEN_344;
  wire [31:0] _GEN_345;
  wire [31:0] _GEN_346;
  wire [31:0] _GEN_347;
  wire [31:0] _GEN_348;
  wire [31:0] _GEN_349;
  wire [31:0] _GEN_350;
  wire [31:0] _GEN_351;
  wire [31:0] _GEN_352;
  wire [31:0] _GEN_353;
  wire [31:0] _GEN_354;
  wire [31:0] _GEN_355;
  wire [31:0] _GEN_356;
  wire [31:0] _GEN_357;
  wire [31:0] _GEN_358;
  wire [31:0] _GEN_359;
  wire [31:0] _GEN_360;
  wire [31:0] _GEN_361;
  wire [31:0] _GEN_362;
  wire [31:0] _GEN_363;
  wire [31:0] _GEN_364;
  wire [31:0] _GEN_365;
  wire [31:0] _GEN_366;
  wire [31:0] _GEN_367;
  wire [31:0] _GEN_368;
  wire [31:0] _GEN_369;
  wire [31:0] _GEN_370;
  wire [31:0] _GEN_371;
  wire [31:0] _GEN_372;
  wire [31:0] _GEN_373;
  wire [1:0] _T_12385;
  wire [1:0] _T_12386;
  wire  _T_12387;
  wire  _T_12388;
  wire  _T_12390;
  wire  _T_12391;
  wire  _T_12393;
  wire  _T_12395;
  reg  _T_12398;
  reg [31:0] _RAND_128;
  reg  _T_12412_0;
  reg [31:0] _RAND_129;
  reg  _T_12433_0;
  reg [31:0] _RAND_130;
  reg [31:0] _T_12514_0_0;
  reg [31:0] _RAND_131;
  reg [31:0] _T_12514_0_1;
  reg [31:0] _RAND_132;
  reg [31:0] _T_12514_0_2;
  reg [31:0] _RAND_133;
  reg [31:0] _T_12514_0_3;
  reg [31:0] _RAND_134;
  reg [31:0] _T_12514_0_4;
  reg [31:0] _RAND_135;
  reg [31:0] _T_12514_0_5;
  reg [31:0] _RAND_136;
  reg [31:0] _T_12514_0_6;
  reg [31:0] _RAND_137;
  reg [31:0] _T_12514_0_7;
  reg [31:0] _RAND_138;
  reg [31:0] _T_12514_0_8;
  reg [31:0] _RAND_139;
  reg [31:0] _T_12514_0_9;
  reg [31:0] _RAND_140;
  reg [31:0] _T_12514_0_10;
  reg [31:0] _RAND_141;
  reg [31:0] _T_12514_0_11;
  reg [31:0] _RAND_142;
  reg [31:0] _T_12514_0_12;
  reg [31:0] _RAND_143;
  reg [31:0] _T_12514_0_13;
  reg [31:0] _RAND_144;
  reg [31:0] _T_12514_0_14;
  reg [31:0] _RAND_145;
  reg [31:0] _T_12514_0_15;
  reg [31:0] _RAND_146;
  reg [31:0] _T_12514_0_16;
  reg [31:0] _RAND_147;
  reg [31:0] _T_12514_0_17;
  reg [31:0] _RAND_148;
  reg [31:0] _T_12514_0_18;
  reg [31:0] _RAND_149;
  reg [31:0] _T_12514_0_19;
  reg [31:0] _RAND_150;
  reg [31:0] _T_12514_0_20;
  reg [31:0] _RAND_151;
  reg [31:0] _T_12514_0_21;
  reg [31:0] _RAND_152;
  reg [31:0] _T_12514_0_22;
  reg [31:0] _RAND_153;
  reg [31:0] _T_12514_0_23;
  reg [31:0] _RAND_154;
  reg [31:0] _T_12514_0_24;
  reg [31:0] _RAND_155;
  reg [31:0] _T_12514_0_25;
  reg [31:0] _RAND_156;
  reg [31:0] _T_12514_0_26;
  reg [31:0] _RAND_157;
  reg [31:0] _T_12514_0_27;
  reg [31:0] _RAND_158;
  reg [31:0] _T_12514_0_28;
  reg [31:0] _RAND_159;
  reg [31:0] _T_12514_0_29;
  reg [31:0] _RAND_160;
  reg [31:0] _T_12514_0_30;
  reg [31:0] _RAND_161;
  reg [31:0] _T_12514_0_31;
  reg [31:0] _RAND_162;
  reg [4:0] _T_12733_0;
  reg [31:0] _RAND_163;
  reg  _T_12754_0;
  reg [31:0] _RAND_164;
  reg  _T_12764;
  reg [31:0] _RAND_165;
  reg  _T_12767;
  reg [31:0] _RAND_166;
  reg  _T_12770;
  reg [31:0] _RAND_167;
  wire  _T_12774;
  wire  _T_12776;
  wire [1:0] _T_12778;
  wire  _T_12779;
  wire  _GEN_374;
  wire  _T_12786;
  wire  _T_12792;
  wire  _T_12793;
  wire  _T_12795;
  wire  _T_12800;
  wire  _T_12807;
  wire  _T_12808;
  wire  _GEN_375;
  wire  _T_12820;
  wire [1:0] _T_12831;
  wire  _T_12832;
  wire  _GEN_377;
  wire  _GEN_378;
  wire  _GEN_379;
  wire  _GEN_380;
  wire  _GEN_382;
  wire  _GEN_383;
  wire  _T_12834;
  wire [5:0] _T_12840;
  wire [4:0] _T_12841;
  wire  _GEN_384;
  wire  _GEN_385;
  wire  _GEN_386;
  wire [4:0] _GEN_387;
  wire  _GEN_388;
  wire  _GEN_389;
  wire  _GEN_390;
  wire [4:0] _GEN_391;
  wire  _T_12842;
  wire [1:0] _T_12847;
  wire  _T_12848;
  wire  _T_12849;
  wire  _T_12851;
  wire [31:0] _T_12955;
  wire [31:0] _GEN_392;
  wire [31:0] _T_13061;
  wire [31:0] _GEN_393;
  wire [31:0] _T_13167;
  wire [31:0] _GEN_394;
  wire [31:0] _T_13273;
  wire [31:0] _GEN_395;
  wire [31:0] _T_13379;
  wire [31:0] _GEN_396;
  wire [31:0] _T_13485;
  wire [31:0] _GEN_397;
  wire [31:0] _T_13591;
  wire [31:0] _GEN_398;
  wire [31:0] _T_13697;
  wire [31:0] _GEN_399;
  wire [31:0] _T_13803;
  wire [31:0] _GEN_400;
  wire [31:0] _T_13909;
  wire [31:0] _GEN_401;
  wire [31:0] _T_14015;
  wire [31:0] _GEN_402;
  wire [31:0] _T_14121;
  wire [31:0] _GEN_403;
  wire [31:0] _T_14227;
  wire [31:0] _GEN_404;
  wire [31:0] _T_14333;
  wire [31:0] _GEN_405;
  wire [31:0] _T_14439;
  wire [31:0] _GEN_406;
  wire [31:0] _T_14545;
  wire [31:0] _GEN_407;
  wire [31:0] _GEN_408;
  wire [31:0] _GEN_409;
  wire [31:0] _GEN_410;
  wire [31:0] _GEN_411;
  wire [31:0] _GEN_412;
  wire [31:0] _GEN_413;
  wire [31:0] _GEN_414;
  wire [31:0] _GEN_415;
  wire [31:0] _GEN_416;
  wire [31:0] _GEN_417;
  wire [31:0] _GEN_418;
  wire [31:0] _GEN_419;
  wire [31:0] _GEN_420;
  wire [31:0] _GEN_421;
  wire [31:0] _GEN_422;
  wire [31:0] _GEN_423;
  wire  _GEN_424;
  wire [31:0] _GEN_425;
  wire [31:0] _GEN_426;
  wire [31:0] _GEN_427;
  wire [31:0] _GEN_428;
  wire [31:0] _GEN_429;
  wire [31:0] _GEN_430;
  wire [31:0] _GEN_431;
  wire [31:0] _GEN_432;
  wire [31:0] _GEN_433;
  wire [31:0] _GEN_434;
  wire [31:0] _GEN_435;
  wire [31:0] _GEN_436;
  wire [31:0] _GEN_437;
  wire [31:0] _GEN_438;
  wire [31:0] _GEN_439;
  wire [31:0] _GEN_440;
  wire [31:0] _GEN_441;
  wire [31:0] _GEN_442;
  wire [31:0] _GEN_443;
  wire [31:0] _GEN_444;
  wire [31:0] _GEN_445;
  wire [31:0] _GEN_446;
  wire [31:0] _GEN_447;
  wire [31:0] _GEN_448;
  wire [31:0] _GEN_449;
  wire [31:0] _GEN_450;
  wire [31:0] _GEN_451;
  wire [31:0] _GEN_452;
  wire [31:0] _GEN_453;
  wire [31:0] _GEN_454;
  wire [31:0] _GEN_455;
  wire [31:0] _GEN_456;
  wire  _T_16242;
  wire  _T_16245;
  wire  _T_16255;
  wire  _T_16256;
  wire  _T_16262;
  wire  _T_16263;
  wire  _T_16264;
  wire  _GEN_457;
  wire  _GEN_458;
  wire  _T_16276;
  wire  _T_16278;
  wire [1:0] _T_16281;
  wire  _T_16282;
  wire  _T_16283;
  wire [1:0] _T_16286;
  wire  _T_16287;
  wire  _GEN_459;
  wire  _GEN_460;
  wire  _GEN_461;
  wire  _GEN_462;
  wire  _GEN_463;
  wire  _GEN_464;
  wire  _T_16298;
  wire [31:0] _GEN_3;
  wire [31:0] _GEN_465;
  wire [31:0] _GEN_466;
  wire [31:0] _GEN_467;
  wire [31:0] _GEN_468;
  wire [31:0] _GEN_469;
  wire [31:0] _GEN_470;
  wire [31:0] _GEN_471;
  wire [31:0] _GEN_472;
  wire [31:0] _GEN_473;
  wire [31:0] _GEN_474;
  wire [31:0] _GEN_475;
  wire [31:0] _GEN_476;
  wire [31:0] _GEN_477;
  wire [31:0] _GEN_478;
  wire [31:0] _GEN_479;
  wire [31:0] _GEN_480;
  wire [31:0] _GEN_481;
  wire [31:0] _GEN_482;
  wire [31:0] _GEN_483;
  wire [31:0] _GEN_484;
  wire [31:0] _GEN_485;
  wire [31:0] _GEN_486;
  wire [31:0] _GEN_487;
  wire [31:0] _GEN_488;
  wire [31:0] _GEN_489;
  wire [31:0] _GEN_490;
  wire [31:0] _GEN_491;
  wire [31:0] _GEN_492;
  wire [31:0] _GEN_493;
  wire [31:0] _GEN_494;
  wire [31:0] _GEN_495;
  wire [1:0] _T_16305;
  wire [1:0] _T_16306;
  wire  _T_16307;
  wire  _T_16308;
  wire  _T_16310;
  wire  _T_16311;
  wire  _T_16313;
  wire  _T_16315;
  reg  _T_16318;
  reg [31:0] _RAND_168;
  wire [1:0] _T_16322;
  wire  _T_16323;
  wire  _GEN_496;
  reg  _T_16337_0;
  reg [31:0] _RAND_169;
  wire  _T_16346;
  reg [31:0] _T_16350_0;
  reg [31:0] _RAND_170;
  reg [31:0] _T_16427_0_0;
  reg [31:0] _RAND_171;
  reg [31:0] _T_16427_0_1;
  reg [31:0] _RAND_172;
  reg [31:0] _T_16427_0_2;
  reg [31:0] _RAND_173;
  reg [31:0] _T_16427_0_3;
  reg [31:0] _RAND_174;
  reg [31:0] _T_16427_0_4;
  reg [31:0] _RAND_175;
  reg [31:0] _T_16427_0_5;
  reg [31:0] _RAND_176;
  reg [31:0] _T_16427_0_6;
  reg [31:0] _RAND_177;
  reg [31:0] _T_16427_0_7;
  reg [31:0] _RAND_178;
  reg [31:0] _T_16427_0_8;
  reg [31:0] _RAND_179;
  reg [31:0] _T_16427_0_9;
  reg [31:0] _RAND_180;
  reg [31:0] _T_16427_0_10;
  reg [31:0] _RAND_181;
  reg [31:0] _T_16427_0_11;
  reg [31:0] _RAND_182;
  reg [31:0] _T_16427_0_12;
  reg [31:0] _RAND_183;
  reg [31:0] _T_16427_0_13;
  reg [31:0] _RAND_184;
  reg [31:0] _T_16427_0_14;
  reg [31:0] _RAND_185;
  reg [31:0] _T_16427_0_15;
  reg [31:0] _RAND_186;
  reg [31:0] _T_16427_0_16;
  reg [31:0] _RAND_187;
  reg [31:0] _T_16427_0_17;
  reg [31:0] _RAND_188;
  reg [31:0] _T_16427_0_18;
  reg [31:0] _RAND_189;
  reg [31:0] _T_16427_0_19;
  reg [31:0] _RAND_190;
  reg [31:0] _T_16427_0_20;
  reg [31:0] _RAND_191;
  reg [31:0] _T_16427_0_21;
  reg [31:0] _RAND_192;
  reg [31:0] _T_16427_0_22;
  reg [31:0] _RAND_193;
  reg [31:0] _T_16427_0_23;
  reg [31:0] _RAND_194;
  reg [31:0] _T_16427_0_24;
  reg [31:0] _RAND_195;
  reg [31:0] _T_16427_0_25;
  reg [31:0] _RAND_196;
  reg [31:0] _T_16427_0_26;
  reg [31:0] _RAND_197;
  reg [31:0] _T_16427_0_27;
  reg [31:0] _RAND_198;
  reg [31:0] _T_16427_0_28;
  reg [31:0] _RAND_199;
  reg [31:0] _T_16427_0_29;
  reg [31:0] _RAND_200;
  reg [31:0] _T_16427_0_30;
  reg [31:0] _RAND_201;
  reg [31:0] _T_16427_0_31;
  reg [31:0] _RAND_202;
  reg  _T_16646_0;
  reg [31:0] _RAND_203;
  reg  _T_16656;
  reg [31:0] _RAND_204;
  reg  _T_16659;
  reg [31:0] _RAND_205;
  reg  _T_16662;
  reg [31:0] _RAND_206;
  reg  _T_16665;
  reg [31:0] _RAND_207;
  reg  _T_16668;
  reg [31:0] _RAND_208;
  wire  _T_16670;
  wire  _T_16672;
  wire  _T_16673;
  wire  _GEN_497;
  wire  _T_16677;
  wire  _T_16679;
  wire  _T_16680;
  wire  _GEN_498;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_499;
  wire [31:0] _GEN_500;
  wire [31:0] _GEN_501;
  wire [31:0] _GEN_502;
  wire [31:0] _GEN_503;
  wire [31:0] _GEN_504;
  wire [31:0] _GEN_505;
  wire [31:0] _GEN_506;
  wire [31:0] _GEN_507;
  wire [31:0] _GEN_508;
  wire [31:0] _GEN_509;
  wire [31:0] _GEN_510;
  wire [31:0] _GEN_511;
  wire [31:0] _GEN_512;
  wire [31:0] _GEN_513;
  wire [31:0] _GEN_514;
  wire [31:0] _GEN_515;
  wire [31:0] _GEN_516;
  wire [31:0] _GEN_517;
  wire [31:0] _GEN_518;
  wire [31:0] _GEN_519;
  wire [31:0] _GEN_520;
  wire [31:0] _GEN_521;
  wire [31:0] _GEN_522;
  wire [31:0] _GEN_523;
  wire [31:0] _GEN_524;
  wire [31:0] _GEN_525;
  wire [31:0] _GEN_526;
  wire [31:0] _GEN_527;
  wire [31:0] _GEN_528;
  wire [31:0] _GEN_529;
  wire [31:0] _GEN_530;
  wire [31:0] _GEN_531;
  wire [31:0] _GEN_532;
  wire [31:0] _GEN_533;
  wire [31:0] _GEN_534;
  wire [31:0] _GEN_535;
  wire [31:0] _GEN_536;
  wire [31:0] _GEN_537;
  wire [31:0] _GEN_538;
  wire [31:0] _GEN_539;
  wire [31:0] _GEN_540;
  wire [31:0] _GEN_541;
  wire [31:0] _GEN_542;
  wire [31:0] _GEN_543;
  wire [31:0] _GEN_544;
  wire [31:0] _GEN_545;
  wire [31:0] _GEN_546;
  wire [31:0] _GEN_547;
  wire [31:0] _GEN_548;
  wire [31:0] _GEN_549;
  wire [31:0] _GEN_550;
  wire [31:0] _GEN_551;
  wire [31:0] _GEN_552;
  wire [31:0] _GEN_553;
  wire [31:0] _GEN_554;
  wire [31:0] _GEN_555;
  wire [31:0] _GEN_556;
  wire [31:0] _GEN_557;
  wire [31:0] _GEN_558;
  wire [31:0] _GEN_559;
  wire [31:0] _GEN_560;
  wire [31:0] _GEN_561;
  wire [31:0] _GEN_562;
  wire  _T_16686;
  wire  _T_16689;
  wire  _T_16695;
  wire  _GEN_563;
  wire [31:0] _GEN_564;
  wire  _T_16704;
  wire  _T_16705;
  wire [63:0] _T_16810;
  wire [63:0] _T_16811;
  wire [127:0] _T_16812;
  wire [63:0] _T_16813;
  wire [63:0] _T_16814;
  wire [127:0] _T_16815;
  wire [255:0] _T_16816;
  wire [63:0] _T_16817;
  wire [63:0] _T_16818;
  wire [127:0] _T_16819;
  wire [63:0] _T_16820;
  wire [63:0] _T_16821;
  wire [127:0] _T_16822;
  wire [255:0] _T_16823;
  wire [511:0] _T_16824;
  wire [63:0] _T_16825;
  wire [63:0] _T_16826;
  wire [127:0] _T_16827;
  wire [63:0] _T_16828;
  wire [63:0] _T_16829;
  wire [127:0] _T_16830;
  wire [255:0] _T_16831;
  wire [63:0] _T_16832;
  wire [63:0] _T_16833;
  wire [127:0] _T_16834;
  wire [63:0] _T_16835;
  wire [63:0] _T_16836;
  wire [127:0] _T_16837;
  wire [255:0] _T_16838;
  wire [511:0] _T_16839;
  wire [1023:0] _T_16840;
  wire [511:0] _T_16841;
  wire [511:0] _T_16844;
  wire [511:0] _T_16845;
  wire  _T_16852;
  wire  _T_16859;
  wire  _T_16860;
  wire  _T_16862;
  wire [1:0] _T_16865;
  wire  _T_16866;
  wire  _GEN_565;
  wire  _GEN_566;
  wire  _GEN_567;
  wire  _GEN_568;
  wire  _T_16867;
  wire [1:0] _T_16872;
  wire  _T_16873;
  wire  _T_16874;
  wire  _GEN_569;
  wire  _T_16878;
  wire  _T_16885;
  wire  _T_16886;
  wire  _T_16887;
  wire  _T_16888;
  wire  _T_16890;
  wire  _T_16892;
  wire [1:0] _T_16895;
  wire  _T_16896;
  wire  _T_16897;
  wire [1:0] _T_16906;
  wire  _T_16907;
  wire  _GEN_570;
  wire  _GEN_571;
  wire  _GEN_572;
  wire  _GEN_573;
  wire  _GEN_574;
  wire  _GEN_575;
  wire  _GEN_576;
  wire  _GEN_577;
  wire  _GEN_578;
  wire  _GEN_579;
  wire  _GEN_580;
  wire  _GEN_581;
  wire  _GEN_582;
  wire  _GEN_583;
  wire  _GEN_584;
  wire  _GEN_585;
  wire  _T_16923;
  reg  _T_16926;
  reg [31:0] _RAND_209;
  wire [1:0] _T_16930;
  wire  _T_16931;
  wire  _GEN_586;
  reg  _T_16945_0;
  reg [31:0] _RAND_210;
  wire  _T_16954;
  reg [31:0] _T_16958_0;
  reg [31:0] _RAND_211;
  reg [31:0] _T_17035_0_0;
  reg [31:0] _RAND_212;
  reg [31:0] _T_17035_0_1;
  reg [31:0] _RAND_213;
  reg [31:0] _T_17035_0_2;
  reg [31:0] _RAND_214;
  reg [31:0] _T_17035_0_3;
  reg [31:0] _RAND_215;
  reg [31:0] _T_17035_0_4;
  reg [31:0] _RAND_216;
  reg [31:0] _T_17035_0_5;
  reg [31:0] _RAND_217;
  reg [31:0] _T_17035_0_6;
  reg [31:0] _RAND_218;
  reg [31:0] _T_17035_0_7;
  reg [31:0] _RAND_219;
  reg [31:0] _T_17035_0_8;
  reg [31:0] _RAND_220;
  reg [31:0] _T_17035_0_9;
  reg [31:0] _RAND_221;
  reg [31:0] _T_17035_0_10;
  reg [31:0] _RAND_222;
  reg [31:0] _T_17035_0_11;
  reg [31:0] _RAND_223;
  reg [31:0] _T_17035_0_12;
  reg [31:0] _RAND_224;
  reg [31:0] _T_17035_0_13;
  reg [31:0] _RAND_225;
  reg [31:0] _T_17035_0_14;
  reg [31:0] _RAND_226;
  reg [31:0] _T_17035_0_15;
  reg [31:0] _RAND_227;
  reg [31:0] _T_17035_0_16;
  reg [31:0] _RAND_228;
  reg [31:0] _T_17035_0_17;
  reg [31:0] _RAND_229;
  reg [31:0] _T_17035_0_18;
  reg [31:0] _RAND_230;
  reg [31:0] _T_17035_0_19;
  reg [31:0] _RAND_231;
  reg [31:0] _T_17035_0_20;
  reg [31:0] _RAND_232;
  reg [31:0] _T_17035_0_21;
  reg [31:0] _RAND_233;
  reg [31:0] _T_17035_0_22;
  reg [31:0] _RAND_234;
  reg [31:0] _T_17035_0_23;
  reg [31:0] _RAND_235;
  reg [31:0] _T_17035_0_24;
  reg [31:0] _RAND_236;
  reg [31:0] _T_17035_0_25;
  reg [31:0] _RAND_237;
  reg [31:0] _T_17035_0_26;
  reg [31:0] _RAND_238;
  reg [31:0] _T_17035_0_27;
  reg [31:0] _RAND_239;
  reg [31:0] _T_17035_0_28;
  reg [31:0] _RAND_240;
  reg [31:0] _T_17035_0_29;
  reg [31:0] _RAND_241;
  reg [31:0] _T_17035_0_30;
  reg [31:0] _RAND_242;
  reg [31:0] _T_17035_0_31;
  reg [31:0] _RAND_243;
  reg  _T_17254_0;
  reg [31:0] _RAND_244;
  reg  _T_17264;
  reg [31:0] _RAND_245;
  reg  _T_17267;
  reg [31:0] _RAND_246;
  reg  _T_17270;
  reg [31:0] _RAND_247;
  reg  _T_17273;
  reg [31:0] _RAND_248;
  reg  _T_17276;
  reg [31:0] _RAND_249;
  wire  _T_17278;
  wire  _T_17280;
  wire  _T_17281;
  wire  _GEN_587;
  wire  _T_17285;
  wire  _T_17287;
  wire  _T_17288;
  wire  _GEN_588;
  wire [31:0] _GEN_5;
  wire [31:0] _GEN_589;
  wire [31:0] _GEN_590;
  wire [31:0] _GEN_591;
  wire [31:0] _GEN_592;
  wire [31:0] _GEN_593;
  wire [31:0] _GEN_594;
  wire [31:0] _GEN_595;
  wire [31:0] _GEN_596;
  wire [31:0] _GEN_597;
  wire [31:0] _GEN_598;
  wire [31:0] _GEN_599;
  wire [31:0] _GEN_600;
  wire [31:0] _GEN_601;
  wire [31:0] _GEN_602;
  wire [31:0] _GEN_603;
  wire [31:0] _GEN_604;
  wire [31:0] _GEN_605;
  wire [31:0] _GEN_606;
  wire [31:0] _GEN_607;
  wire [31:0] _GEN_608;
  wire [31:0] _GEN_609;
  wire [31:0] _GEN_610;
  wire [31:0] _GEN_611;
  wire [31:0] _GEN_612;
  wire [31:0] _GEN_613;
  wire [31:0] _GEN_614;
  wire [31:0] _GEN_615;
  wire [31:0] _GEN_616;
  wire [31:0] _GEN_617;
  wire [31:0] _GEN_618;
  wire [31:0] _GEN_619;
  wire [31:0] _GEN_620;
  wire [31:0] _GEN_621;
  wire [31:0] _GEN_622;
  wire [31:0] _GEN_623;
  wire [31:0] _GEN_624;
  wire [31:0] _GEN_625;
  wire [31:0] _GEN_626;
  wire [31:0] _GEN_627;
  wire [31:0] _GEN_628;
  wire [31:0] _GEN_629;
  wire [31:0] _GEN_630;
  wire [31:0] _GEN_631;
  wire [31:0] _GEN_632;
  wire [31:0] _GEN_633;
  wire [31:0] _GEN_634;
  wire [31:0] _GEN_635;
  wire [31:0] _GEN_636;
  wire [31:0] _GEN_637;
  wire [31:0] _GEN_638;
  wire [31:0] _GEN_639;
  wire [31:0] _GEN_640;
  wire [31:0] _GEN_641;
  wire [31:0] _GEN_642;
  wire [31:0] _GEN_643;
  wire [31:0] _GEN_644;
  wire [31:0] _GEN_645;
  wire [31:0] _GEN_646;
  wire [31:0] _GEN_647;
  wire [31:0] _GEN_648;
  wire [31:0] _GEN_649;
  wire [31:0] _GEN_650;
  wire [31:0] _GEN_651;
  wire [31:0] _GEN_652;
  wire  _T_17294;
  wire  _T_17297;
  wire  _T_17303;
  wire  _GEN_653;
  wire [31:0] _GEN_654;
  wire  _T_17312;
  wire  _T_17313;
  wire [63:0] _T_17418;
  wire [63:0] _T_17419;
  wire [127:0] _T_17420;
  wire [63:0] _T_17421;
  wire [63:0] _T_17422;
  wire [127:0] _T_17423;
  wire [255:0] _T_17424;
  wire [63:0] _T_17425;
  wire [63:0] _T_17426;
  wire [127:0] _T_17427;
  wire [63:0] _T_17428;
  wire [63:0] _T_17429;
  wire [127:0] _T_17430;
  wire [255:0] _T_17431;
  wire [511:0] _T_17432;
  wire [63:0] _T_17433;
  wire [63:0] _T_17434;
  wire [127:0] _T_17435;
  wire [63:0] _T_17436;
  wire [63:0] _T_17437;
  wire [127:0] _T_17438;
  wire [255:0] _T_17439;
  wire [63:0] _T_17440;
  wire [63:0] _T_17441;
  wire [127:0] _T_17442;
  wire [63:0] _T_17443;
  wire [63:0] _T_17444;
  wire [127:0] _T_17445;
  wire [255:0] _T_17446;
  wire [511:0] _T_17447;
  wire [1023:0] _T_17448;
  wire [511:0] _T_17449;
  wire [511:0] _T_17452;
  wire [511:0] _T_17453;
  wire  _T_17460;
  wire  _T_17467;
  wire  _T_17468;
  wire  _T_17470;
  wire [1:0] _T_17473;
  wire  _T_17474;
  wire  _GEN_655;
  wire  _GEN_656;
  wire  _GEN_657;
  wire  _GEN_658;
  wire  _T_17475;
  wire [1:0] _T_17480;
  wire  _T_17481;
  wire  _T_17482;
  wire  _GEN_659;
  wire  _T_17486;
  wire  _T_17493;
  wire  _T_17494;
  wire  _T_17495;
  wire  _T_17496;
  wire  _T_17498;
  wire  _T_17500;
  wire [1:0] _T_17503;
  wire  _T_17504;
  wire  _T_17505;
  wire [1:0] _T_17514;
  wire  _T_17515;
  wire  _GEN_660;
  wire  _GEN_661;
  wire  _GEN_662;
  wire  _GEN_663;
  wire  _GEN_664;
  wire  _GEN_665;
  wire  _GEN_666;
  wire  _GEN_667;
  wire  _GEN_668;
  wire  _GEN_669;
  wire  _GEN_670;
  wire  _GEN_671;
  wire  _GEN_672;
  wire  _GEN_673;
  wire  _GEN_674;
  wire  _GEN_675;
  wire  _T_17531;
  reg  _T_17534;
  reg [31:0] _RAND_250;
  wire [1:0] _T_17538;
  wire  _T_17539;
  wire  _GEN_676;
  reg  _T_17553_0;
  reg [31:0] _RAND_251;
  wire  _T_17562;
  reg [31:0] _T_17566_0;
  reg [31:0] _RAND_252;
  reg [31:0] _T_17643_0_0;
  reg [31:0] _RAND_253;
  reg [31:0] _T_17643_0_1;
  reg [31:0] _RAND_254;
  reg [31:0] _T_17643_0_2;
  reg [31:0] _RAND_255;
  reg [31:0] _T_17643_0_3;
  reg [31:0] _RAND_256;
  reg [31:0] _T_17643_0_4;
  reg [31:0] _RAND_257;
  reg [31:0] _T_17643_0_5;
  reg [31:0] _RAND_258;
  reg [31:0] _T_17643_0_6;
  reg [31:0] _RAND_259;
  reg [31:0] _T_17643_0_7;
  reg [31:0] _RAND_260;
  reg [31:0] _T_17643_0_8;
  reg [31:0] _RAND_261;
  reg [31:0] _T_17643_0_9;
  reg [31:0] _RAND_262;
  reg [31:0] _T_17643_0_10;
  reg [31:0] _RAND_263;
  reg [31:0] _T_17643_0_11;
  reg [31:0] _RAND_264;
  reg [31:0] _T_17643_0_12;
  reg [31:0] _RAND_265;
  reg [31:0] _T_17643_0_13;
  reg [31:0] _RAND_266;
  reg [31:0] _T_17643_0_14;
  reg [31:0] _RAND_267;
  reg [31:0] _T_17643_0_15;
  reg [31:0] _RAND_268;
  reg [31:0] _T_17643_0_16;
  reg [31:0] _RAND_269;
  reg [31:0] _T_17643_0_17;
  reg [31:0] _RAND_270;
  reg [31:0] _T_17643_0_18;
  reg [31:0] _RAND_271;
  reg [31:0] _T_17643_0_19;
  reg [31:0] _RAND_272;
  reg [31:0] _T_17643_0_20;
  reg [31:0] _RAND_273;
  reg [31:0] _T_17643_0_21;
  reg [31:0] _RAND_274;
  reg [31:0] _T_17643_0_22;
  reg [31:0] _RAND_275;
  reg [31:0] _T_17643_0_23;
  reg [31:0] _RAND_276;
  reg [31:0] _T_17643_0_24;
  reg [31:0] _RAND_277;
  reg [31:0] _T_17643_0_25;
  reg [31:0] _RAND_278;
  reg [31:0] _T_17643_0_26;
  reg [31:0] _RAND_279;
  reg [31:0] _T_17643_0_27;
  reg [31:0] _RAND_280;
  reg [31:0] _T_17643_0_28;
  reg [31:0] _RAND_281;
  reg [31:0] _T_17643_0_29;
  reg [31:0] _RAND_282;
  reg [31:0] _T_17643_0_30;
  reg [31:0] _RAND_283;
  reg [31:0] _T_17643_0_31;
  reg [31:0] _RAND_284;
  reg  _T_17862_0;
  reg [31:0] _RAND_285;
  reg  _T_17872;
  reg [31:0] _RAND_286;
  reg  _T_17875;
  reg [31:0] _RAND_287;
  reg  _T_17878;
  reg [31:0] _RAND_288;
  reg  _T_17881;
  reg [31:0] _RAND_289;
  reg  _T_17884;
  reg [31:0] _RAND_290;
  wire  _T_17886;
  wire  _T_17888;
  wire  _T_17889;
  wire  _GEN_677;
  wire  _T_17893;
  wire  _T_17895;
  wire  _T_17896;
  wire  _GEN_678;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_679;
  wire [31:0] _GEN_680;
  wire [31:0] _GEN_681;
  wire [31:0] _GEN_682;
  wire [31:0] _GEN_683;
  wire [31:0] _GEN_684;
  wire [31:0] _GEN_685;
  wire [31:0] _GEN_686;
  wire [31:0] _GEN_687;
  wire [31:0] _GEN_688;
  wire [31:0] _GEN_689;
  wire [31:0] _GEN_690;
  wire [31:0] _GEN_691;
  wire [31:0] _GEN_692;
  wire [31:0] _GEN_693;
  wire [31:0] _GEN_694;
  wire [31:0] _GEN_695;
  wire [31:0] _GEN_696;
  wire [31:0] _GEN_697;
  wire [31:0] _GEN_698;
  wire [31:0] _GEN_699;
  wire [31:0] _GEN_700;
  wire [31:0] _GEN_701;
  wire [31:0] _GEN_702;
  wire [31:0] _GEN_703;
  wire [31:0] _GEN_704;
  wire [31:0] _GEN_705;
  wire [31:0] _GEN_706;
  wire [31:0] _GEN_707;
  wire [31:0] _GEN_708;
  wire [31:0] _GEN_709;
  wire [31:0] _GEN_710;
  wire [31:0] _GEN_711;
  wire [31:0] _GEN_712;
  wire [31:0] _GEN_713;
  wire [31:0] _GEN_714;
  wire [31:0] _GEN_715;
  wire [31:0] _GEN_716;
  wire [31:0] _GEN_717;
  wire [31:0] _GEN_718;
  wire [31:0] _GEN_719;
  wire [31:0] _GEN_720;
  wire [31:0] _GEN_721;
  wire [31:0] _GEN_722;
  wire [31:0] _GEN_723;
  wire [31:0] _GEN_724;
  wire [31:0] _GEN_725;
  wire [31:0] _GEN_726;
  wire [31:0] _GEN_727;
  wire [31:0] _GEN_728;
  wire [31:0] _GEN_729;
  wire [31:0] _GEN_730;
  wire [31:0] _GEN_731;
  wire [31:0] _GEN_732;
  wire [31:0] _GEN_733;
  wire [31:0] _GEN_734;
  wire [31:0] _GEN_735;
  wire [31:0] _GEN_736;
  wire [31:0] _GEN_737;
  wire [31:0] _GEN_738;
  wire [31:0] _GEN_739;
  wire [31:0] _GEN_740;
  wire [31:0] _GEN_741;
  wire [31:0] _GEN_742;
  wire  _T_17902;
  wire  _T_17905;
  wire  _T_17911;
  wire  _GEN_743;
  wire [31:0] _GEN_744;
  wire  _T_17920;
  wire  _T_17921;
  wire [63:0] _T_18026;
  wire [63:0] _T_18027;
  wire [127:0] _T_18028;
  wire [63:0] _T_18029;
  wire [63:0] _T_18030;
  wire [127:0] _T_18031;
  wire [255:0] _T_18032;
  wire [63:0] _T_18033;
  wire [63:0] _T_18034;
  wire [127:0] _T_18035;
  wire [63:0] _T_18036;
  wire [63:0] _T_18037;
  wire [127:0] _T_18038;
  wire [255:0] _T_18039;
  wire [511:0] _T_18040;
  wire [63:0] _T_18041;
  wire [63:0] _T_18042;
  wire [127:0] _T_18043;
  wire [63:0] _T_18044;
  wire [63:0] _T_18045;
  wire [127:0] _T_18046;
  wire [255:0] _T_18047;
  wire [63:0] _T_18048;
  wire [63:0] _T_18049;
  wire [127:0] _T_18050;
  wire [63:0] _T_18051;
  wire [63:0] _T_18052;
  wire [127:0] _T_18053;
  wire [255:0] _T_18054;
  wire [511:0] _T_18055;
  wire [1023:0] _T_18056;
  wire [511:0] _T_18057;
  wire [511:0] _T_18060;
  wire [511:0] _T_18061;
  wire  _T_18068;
  wire  _T_18075;
  wire  _T_18076;
  wire  _T_18078;
  wire [1:0] _T_18081;
  wire  _T_18082;
  wire  _GEN_745;
  wire  _GEN_746;
  wire  _GEN_747;
  wire  _GEN_748;
  wire  _T_18083;
  wire [1:0] _T_18088;
  wire  _T_18089;
  wire  _T_18090;
  wire  _GEN_749;
  wire  _T_18094;
  wire  _T_18101;
  wire  _T_18102;
  wire  _T_18103;
  wire  _T_18104;
  wire  _T_18106;
  wire  _T_18108;
  wire [1:0] _T_18111;
  wire  _T_18112;
  wire  _T_18113;
  wire [1:0] _T_18122;
  wire  _T_18123;
  wire  _GEN_750;
  wire  _GEN_751;
  wire  _GEN_752;
  wire  _GEN_753;
  wire  _GEN_754;
  wire  _GEN_755;
  wire  _GEN_756;
  wire  _GEN_757;
  wire  _GEN_758;
  wire  _GEN_759;
  wire  _GEN_760;
  wire  _GEN_761;
  wire  _GEN_762;
  wire  _GEN_763;
  wire  _GEN_764;
  wire  _GEN_765;
  wire  _T_18139;
  reg  _T_18142;
  reg [31:0] _RAND_291;
  wire [1:0] _T_18146;
  wire  _T_18147;
  wire  _GEN_766;
  reg  _T_18161_0;
  reg [31:0] _RAND_292;
  wire  _T_18170;
  reg [31:0] _T_18174_0;
  reg [31:0] _RAND_293;
  reg [31:0] _T_18251_0_0;
  reg [31:0] _RAND_294;
  reg [31:0] _T_18251_0_1;
  reg [31:0] _RAND_295;
  reg [31:0] _T_18251_0_2;
  reg [31:0] _RAND_296;
  reg [31:0] _T_18251_0_3;
  reg [31:0] _RAND_297;
  reg [31:0] _T_18251_0_4;
  reg [31:0] _RAND_298;
  reg [31:0] _T_18251_0_5;
  reg [31:0] _RAND_299;
  reg [31:0] _T_18251_0_6;
  reg [31:0] _RAND_300;
  reg [31:0] _T_18251_0_7;
  reg [31:0] _RAND_301;
  reg [31:0] _T_18251_0_8;
  reg [31:0] _RAND_302;
  reg [31:0] _T_18251_0_9;
  reg [31:0] _RAND_303;
  reg [31:0] _T_18251_0_10;
  reg [31:0] _RAND_304;
  reg [31:0] _T_18251_0_11;
  reg [31:0] _RAND_305;
  reg [31:0] _T_18251_0_12;
  reg [31:0] _RAND_306;
  reg [31:0] _T_18251_0_13;
  reg [31:0] _RAND_307;
  reg [31:0] _T_18251_0_14;
  reg [31:0] _RAND_308;
  reg [31:0] _T_18251_0_15;
  reg [31:0] _RAND_309;
  reg [31:0] _T_18251_0_16;
  reg [31:0] _RAND_310;
  reg [31:0] _T_18251_0_17;
  reg [31:0] _RAND_311;
  reg [31:0] _T_18251_0_18;
  reg [31:0] _RAND_312;
  reg [31:0] _T_18251_0_19;
  reg [31:0] _RAND_313;
  reg [31:0] _T_18251_0_20;
  reg [31:0] _RAND_314;
  reg [31:0] _T_18251_0_21;
  reg [31:0] _RAND_315;
  reg [31:0] _T_18251_0_22;
  reg [31:0] _RAND_316;
  reg [31:0] _T_18251_0_23;
  reg [31:0] _RAND_317;
  reg [31:0] _T_18251_0_24;
  reg [31:0] _RAND_318;
  reg [31:0] _T_18251_0_25;
  reg [31:0] _RAND_319;
  reg [31:0] _T_18251_0_26;
  reg [31:0] _RAND_320;
  reg [31:0] _T_18251_0_27;
  reg [31:0] _RAND_321;
  reg [31:0] _T_18251_0_28;
  reg [31:0] _RAND_322;
  reg [31:0] _T_18251_0_29;
  reg [31:0] _RAND_323;
  reg [31:0] _T_18251_0_30;
  reg [31:0] _RAND_324;
  reg [31:0] _T_18251_0_31;
  reg [31:0] _RAND_325;
  reg  _T_18470_0;
  reg [31:0] _RAND_326;
  reg  _T_18480;
  reg [31:0] _RAND_327;
  reg  _T_18483;
  reg [31:0] _RAND_328;
  reg  _T_18486;
  reg [31:0] _RAND_329;
  reg  _T_18489;
  reg [31:0] _RAND_330;
  reg  _T_18492;
  reg [31:0] _RAND_331;
  wire  _T_18494;
  wire  _T_18496;
  wire  _T_18497;
  wire  _GEN_767;
  wire  _T_18501;
  wire  _T_18503;
  wire  _T_18504;
  wire  _GEN_768;
  wire [31:0] _GEN_7;
  wire [31:0] _GEN_769;
  wire [31:0] _GEN_770;
  wire [31:0] _GEN_771;
  wire [31:0] _GEN_772;
  wire [31:0] _GEN_773;
  wire [31:0] _GEN_774;
  wire [31:0] _GEN_775;
  wire [31:0] _GEN_776;
  wire [31:0] _GEN_777;
  wire [31:0] _GEN_778;
  wire [31:0] _GEN_779;
  wire [31:0] _GEN_780;
  wire [31:0] _GEN_781;
  wire [31:0] _GEN_782;
  wire [31:0] _GEN_783;
  wire [31:0] _GEN_784;
  wire [31:0] _GEN_785;
  wire [31:0] _GEN_786;
  wire [31:0] _GEN_787;
  wire [31:0] _GEN_788;
  wire [31:0] _GEN_789;
  wire [31:0] _GEN_790;
  wire [31:0] _GEN_791;
  wire [31:0] _GEN_792;
  wire [31:0] _GEN_793;
  wire [31:0] _GEN_794;
  wire [31:0] _GEN_795;
  wire [31:0] _GEN_796;
  wire [31:0] _GEN_797;
  wire [31:0] _GEN_798;
  wire [31:0] _GEN_799;
  wire [31:0] _GEN_800;
  wire [31:0] _GEN_801;
  wire [31:0] _GEN_802;
  wire [31:0] _GEN_803;
  wire [31:0] _GEN_804;
  wire [31:0] _GEN_805;
  wire [31:0] _GEN_806;
  wire [31:0] _GEN_807;
  wire [31:0] _GEN_808;
  wire [31:0] _GEN_809;
  wire [31:0] _GEN_810;
  wire [31:0] _GEN_811;
  wire [31:0] _GEN_812;
  wire [31:0] _GEN_813;
  wire [31:0] _GEN_814;
  wire [31:0] _GEN_815;
  wire [31:0] _GEN_816;
  wire [31:0] _GEN_817;
  wire [31:0] _GEN_818;
  wire [31:0] _GEN_819;
  wire [31:0] _GEN_820;
  wire [31:0] _GEN_821;
  wire [31:0] _GEN_822;
  wire [31:0] _GEN_823;
  wire [31:0] _GEN_824;
  wire [31:0] _GEN_825;
  wire [31:0] _GEN_826;
  wire [31:0] _GEN_827;
  wire [31:0] _GEN_828;
  wire [31:0] _GEN_829;
  wire [31:0] _GEN_830;
  wire [31:0] _GEN_831;
  wire [31:0] _GEN_832;
  wire  _T_18510;
  wire  _T_18513;
  wire  _T_18519;
  wire  _GEN_833;
  wire [31:0] _GEN_834;
  wire  _T_18528;
  wire  _T_18529;
  wire [63:0] _T_18634;
  wire [63:0] _T_18635;
  wire [127:0] _T_18636;
  wire [63:0] _T_18637;
  wire [63:0] _T_18638;
  wire [127:0] _T_18639;
  wire [255:0] _T_18640;
  wire [63:0] _T_18641;
  wire [63:0] _T_18642;
  wire [127:0] _T_18643;
  wire [63:0] _T_18644;
  wire [63:0] _T_18645;
  wire [127:0] _T_18646;
  wire [255:0] _T_18647;
  wire [511:0] _T_18648;
  wire [63:0] _T_18649;
  wire [63:0] _T_18650;
  wire [127:0] _T_18651;
  wire [63:0] _T_18652;
  wire [63:0] _T_18653;
  wire [127:0] _T_18654;
  wire [255:0] _T_18655;
  wire [63:0] _T_18656;
  wire [63:0] _T_18657;
  wire [127:0] _T_18658;
  wire [63:0] _T_18659;
  wire [63:0] _T_18660;
  wire [127:0] _T_18661;
  wire [255:0] _T_18662;
  wire [511:0] _T_18663;
  wire [1023:0] _T_18664;
  wire [511:0] _T_18665;
  wire [511:0] _T_18668;
  wire [511:0] _T_18669;
  wire  _T_18676;
  wire  _T_18683;
  wire  _T_18684;
  wire  _T_18686;
  wire [1:0] _T_18689;
  wire  _T_18690;
  wire  _GEN_835;
  wire  _GEN_836;
  wire  _GEN_837;
  wire  _GEN_838;
  wire  _T_18691;
  wire [1:0] _T_18696;
  wire  _T_18697;
  wire  _T_18698;
  wire  _GEN_839;
  wire  _T_18702;
  wire  _T_18709;
  wire  _T_18710;
  wire  _T_18711;
  wire  _T_18712;
  wire  _T_18714;
  wire  _T_18716;
  wire [1:0] _T_18719;
  wire  _T_18720;
  wire  _T_18721;
  wire [1:0] _T_18730;
  wire  _T_18731;
  wire  _GEN_840;
  wire  _GEN_841;
  wire  _GEN_842;
  wire  _GEN_843;
  wire  _GEN_844;
  wire  _GEN_845;
  wire  _GEN_846;
  wire  _GEN_847;
  wire  _GEN_848;
  wire  _GEN_849;
  wire  _GEN_850;
  wire  _GEN_851;
  wire  _GEN_852;
  wire  _GEN_853;
  wire  _GEN_854;
  wire  _GEN_855;
  wire  _T_18747;
  wire  _T_18750;
  wire  _T_18751;
  wire  _T_18752;
  wire  _T_18753;
  wire  _T_18754;
  wire  _T_18755;
  wire  cumFinished;
  assign _T_1014 = _T_638 == 1'h0;
  assign _T_1016 = _T_1014 == 1'h0;
  assign _T_1018 = _T_638 + 1'h1;
  assign _T_1019 = _T_1018[0:0];
  assign _GEN_8 = _T_1016 ? _T_1019 : _T_638;
  assign _T_1026 = _T_1014 & _T_428_0;
  assign _T_1032 = _T_652_0 == 1'h0;
  assign _T_1033 = _T_1026 & _T_1032;
  assign _T_1035 = io_axi_inputMemAddrValids_0 & io_axi_inputMemAddrReadys_0;
  assign _T_1040 = _T_1014 & _T_434_0;
  assign _T_1047 = _T_1040 & _T_1032;
  assign _T_1048 = _T_1035 | _T_1047;
  assign _GEN_9 = io_axi_inputMemAddrValids_0 ? 1'h1 : _T_673_0;
  assign _T_1060 = _T_1004 == 1'h0;
  assign _T_1071 = _T_1004 + 1'h1;
  assign _T_1072 = _T_1071[0:0];
  assign _GEN_11 = _T_1060 ? 1'h0 : _GEN_8;
  assign _GEN_12 = _T_1060 ? 1'h0 : _T_1072;
  assign _GEN_13 = _T_1048 ? 1'h1 : _T_652_0;
  assign _GEN_14 = _T_1048 ? _GEN_9 : _T_673_0;
  assign _GEN_16 = _T_1048 ? _GEN_11 : _GEN_8;
  assign _GEN_17 = _T_1048 ? _GEN_12 : _T_1004;
  assign _T_1074 = _T_973_0 == 5'h1f;
  assign _T_1080 = _T_973_0 + 5'h1;
  assign _T_1081 = _T_1080[4:0];
  assign _GEN_18 = _T_1074 ? 1'h0 : _GEN_13;
  assign _GEN_19 = _T_1074 ? 1'h0 : _GEN_14;
  assign _GEN_20 = _T_1074 ? 1'h0 : _T_994_0;
  assign _GEN_21 = _T_1074 ? 5'h0 : _T_1081;
  assign _GEN_22 = _T_994_0 ? _GEN_18 : _GEN_13;
  assign _GEN_23 = _T_994_0 ? _GEN_19 : _GEN_14;
  assign _GEN_24 = _T_994_0 ? _GEN_20 : _T_994_0;
  assign _GEN_25 = _T_994_0 ? _GEN_21 : _T_973_0;
  assign _T_1082 = io_axi_inputMemBlockReadys_0 & io_axi_inputMemBlockValids_0;
  assign _T_1087 = _T_1010 + 1'h1;
  assign _T_1088 = _T_1087[0:0];
  assign _T_1089 = _T_1010 ? 1'h0 : _T_1088;
  assign _T_1091 = 1'h0 == _T_1010;
  assign _T_1195 = io_axi_inputMemBlocks_0[31:0];
  assign _GEN_26 = _T_1091 ? _T_1195 : _T_754_0_0;
  assign _T_1301 = io_axi_inputMemBlocks_0[63:32];
  assign _GEN_27 = _T_1091 ? _T_1301 : _T_754_0_1;
  assign _T_1407 = io_axi_inputMemBlocks_0[95:64];
  assign _GEN_28 = _T_1091 ? _T_1407 : _T_754_0_2;
  assign _T_1513 = io_axi_inputMemBlocks_0[127:96];
  assign _GEN_29 = _T_1091 ? _T_1513 : _T_754_0_3;
  assign _T_1619 = io_axi_inputMemBlocks_0[159:128];
  assign _GEN_30 = _T_1091 ? _T_1619 : _T_754_0_4;
  assign _T_1725 = io_axi_inputMemBlocks_0[191:160];
  assign _GEN_31 = _T_1091 ? _T_1725 : _T_754_0_5;
  assign _T_1831 = io_axi_inputMemBlocks_0[223:192];
  assign _GEN_32 = _T_1091 ? _T_1831 : _T_754_0_6;
  assign _T_1937 = io_axi_inputMemBlocks_0[255:224];
  assign _GEN_33 = _T_1091 ? _T_1937 : _T_754_0_7;
  assign _T_2043 = io_axi_inputMemBlocks_0[287:256];
  assign _GEN_34 = _T_1091 ? _T_2043 : _T_754_0_8;
  assign _T_2149 = io_axi_inputMemBlocks_0[319:288];
  assign _GEN_35 = _T_1091 ? _T_2149 : _T_754_0_9;
  assign _T_2255 = io_axi_inputMemBlocks_0[351:320];
  assign _GEN_36 = _T_1091 ? _T_2255 : _T_754_0_10;
  assign _T_2361 = io_axi_inputMemBlocks_0[383:352];
  assign _GEN_37 = _T_1091 ? _T_2361 : _T_754_0_11;
  assign _T_2467 = io_axi_inputMemBlocks_0[415:384];
  assign _GEN_38 = _T_1091 ? _T_2467 : _T_754_0_12;
  assign _T_2573 = io_axi_inputMemBlocks_0[447:416];
  assign _GEN_39 = _T_1091 ? _T_2573 : _T_754_0_13;
  assign _T_2679 = io_axi_inputMemBlocks_0[479:448];
  assign _GEN_40 = _T_1091 ? _T_2679 : _T_754_0_14;
  assign _T_2785 = io_axi_inputMemBlocks_0[511:480];
  assign _GEN_41 = _T_1091 ? _T_2785 : _T_754_0_15;
  assign _GEN_42 = _T_1010 ? _T_1195 : _T_754_0_16;
  assign _GEN_43 = _T_1010 ? _T_1301 : _T_754_0_17;
  assign _GEN_44 = _T_1010 ? _T_1407 : _T_754_0_18;
  assign _GEN_45 = _T_1010 ? _T_1513 : _T_754_0_19;
  assign _GEN_46 = _T_1010 ? _T_1619 : _T_754_0_20;
  assign _GEN_47 = _T_1010 ? _T_1725 : _T_754_0_21;
  assign _GEN_48 = _T_1010 ? _T_1831 : _T_754_0_22;
  assign _GEN_49 = _T_1010 ? _T_1937 : _T_754_0_23;
  assign _GEN_50 = _T_1010 ? _T_2043 : _T_754_0_24;
  assign _GEN_51 = _T_1010 ? _T_2149 : _T_754_0_25;
  assign _GEN_52 = _T_1010 ? _T_2255 : _T_754_0_26;
  assign _GEN_53 = _T_1010 ? _T_2361 : _T_754_0_27;
  assign _GEN_54 = _T_1010 ? _T_2467 : _T_754_0_28;
  assign _GEN_55 = _T_1010 ? _T_2573 : _T_754_0_29;
  assign _GEN_56 = _T_1010 ? _T_2679 : _T_754_0_30;
  assign _GEN_57 = _T_1010 ? _T_2785 : _T_754_0_31;
  assign _GEN_58 = _T_1082 ? _T_1089 : _T_1010;
  assign _GEN_59 = _T_1082 ? _GEN_26 : _T_754_0_0;
  assign _GEN_60 = _T_1082 ? _GEN_27 : _T_754_0_1;
  assign _GEN_61 = _T_1082 ? _GEN_28 : _T_754_0_2;
  assign _GEN_62 = _T_1082 ? _GEN_29 : _T_754_0_3;
  assign _GEN_63 = _T_1082 ? _GEN_30 : _T_754_0_4;
  assign _GEN_64 = _T_1082 ? _GEN_31 : _T_754_0_5;
  assign _GEN_65 = _T_1082 ? _GEN_32 : _T_754_0_6;
  assign _GEN_66 = _T_1082 ? _GEN_33 : _T_754_0_7;
  assign _GEN_67 = _T_1082 ? _GEN_34 : _T_754_0_8;
  assign _GEN_68 = _T_1082 ? _GEN_35 : _T_754_0_9;
  assign _GEN_69 = _T_1082 ? _GEN_36 : _T_754_0_10;
  assign _GEN_70 = _T_1082 ? _GEN_37 : _T_754_0_11;
  assign _GEN_71 = _T_1082 ? _GEN_38 : _T_754_0_12;
  assign _GEN_72 = _T_1082 ? _GEN_39 : _T_754_0_13;
  assign _GEN_73 = _T_1082 ? _GEN_40 : _T_754_0_14;
  assign _GEN_74 = _T_1082 ? _GEN_41 : _T_754_0_15;
  assign _GEN_75 = _T_1082 ? _GEN_42 : _T_754_0_16;
  assign _GEN_76 = _T_1082 ? _GEN_43 : _T_754_0_17;
  assign _GEN_77 = _T_1082 ? _GEN_44 : _T_754_0_18;
  assign _GEN_78 = _T_1082 ? _GEN_45 : _T_754_0_19;
  assign _GEN_79 = _T_1082 ? _GEN_46 : _T_754_0_20;
  assign _GEN_80 = _T_1082 ? _GEN_47 : _T_754_0_21;
  assign _GEN_81 = _T_1082 ? _GEN_48 : _T_754_0_22;
  assign _GEN_82 = _T_1082 ? _GEN_49 : _T_754_0_23;
  assign _GEN_83 = _T_1082 ? _GEN_50 : _T_754_0_24;
  assign _GEN_84 = _T_1082 ? _GEN_51 : _T_754_0_25;
  assign _GEN_85 = _T_1082 ? _GEN_52 : _T_754_0_26;
  assign _GEN_86 = _T_1082 ? _GEN_53 : _T_754_0_27;
  assign _GEN_87 = _T_1082 ? _GEN_54 : _T_754_0_28;
  assign _GEN_88 = _T_1082 ? _GEN_55 : _T_754_0_29;
  assign _GEN_89 = _T_1082 ? _GEN_56 : _T_754_0_30;
  assign _GEN_90 = _T_1082 ? _GEN_57 : _T_754_0_31;
  assign _T_4482 = io_axi_inputMemBlockValids_0 & io_axi_inputMemBlockReadys_0;
  assign _T_4485 = _T_4482 & _T_1010;
  assign _T_4495 = _T_673_0 == 1'h0;
  assign _T_4496 = _T_652_0 & _T_4495;
  assign _T_4502 = _T_994_0 == 1'h0;
  assign _T_4503 = _T_4496 & _T_4502;
  assign _T_4504 = _T_4485 | _T_4503;
  assign _GEN_91 = io_axi_inputMemBlockReadys_0 ? 1'h1 : _GEN_24;
  assign _GEN_92 = io_axi_inputMemBlockReadys_0 ? _GEN_22 : 1'h0;
  assign _T_4516 = _T_1007 == 1'h0;
  assign _T_4518 = _T_389 == 1'h0;
  assign _T_4521 = _T_389 + 1'h1;
  assign _T_4522 = _T_4521[0:0];
  assign _T_4523 = _T_4518 ? 1'h0 : _T_4522;
  assign _T_4526 = _T_1007 + 1'h1;
  assign _T_4527 = _T_4526[0:0];
  assign _GEN_93 = _T_4516 ? _T_4523 : _T_389;
  assign _GEN_94 = _T_4516 ? 1'h0 : _T_4527;
  assign _GEN_95 = _T_4504 ? _GEN_91 : _GEN_24;
  assign _GEN_96 = _T_4504 ? _GEN_92 : _GEN_22;
  assign _GEN_97 = _T_4504 ? _GEN_93 : _T_389;
  assign _GEN_98 = _T_4504 ? _GEN_94 : _T_1007;
  assign _T_4538 = _T_673_0 & _T_4502;
  assign _GEN_99 = 5'h1 == _T_973_0 ? _T_754_0_1 : _T_754_0_0;
  assign _GEN_100 = 5'h2 == _T_973_0 ? _T_754_0_2 : _GEN_99;
  assign _GEN_101 = 5'h3 == _T_973_0 ? _T_754_0_3 : _GEN_100;
  assign _GEN_102 = 5'h4 == _T_973_0 ? _T_754_0_4 : _GEN_101;
  assign _GEN_103 = 5'h5 == _T_973_0 ? _T_754_0_5 : _GEN_102;
  assign _GEN_104 = 5'h6 == _T_973_0 ? _T_754_0_6 : _GEN_103;
  assign _GEN_105 = 5'h7 == _T_973_0 ? _T_754_0_7 : _GEN_104;
  assign _GEN_106 = 5'h8 == _T_973_0 ? _T_754_0_8 : _GEN_105;
  assign _GEN_107 = 5'h9 == _T_973_0 ? _T_754_0_9 : _GEN_106;
  assign _GEN_108 = 5'ha == _T_973_0 ? _T_754_0_10 : _GEN_107;
  assign _GEN_109 = 5'hb == _T_973_0 ? _T_754_0_11 : _GEN_108;
  assign _GEN_110 = 5'hc == _T_973_0 ? _T_754_0_12 : _GEN_109;
  assign _GEN_111 = 5'hd == _T_973_0 ? _T_754_0_13 : _GEN_110;
  assign _GEN_112 = 5'he == _T_973_0 ? _T_754_0_14 : _GEN_111;
  assign _GEN_113 = 5'hf == _T_973_0 ? _T_754_0_15 : _GEN_112;
  assign _GEN_114 = 5'h10 == _T_973_0 ? _T_754_0_16 : _GEN_113;
  assign _GEN_115 = 5'h11 == _T_973_0 ? _T_754_0_17 : _GEN_114;
  assign _GEN_116 = 5'h12 == _T_973_0 ? _T_754_0_18 : _GEN_115;
  assign _GEN_117 = 5'h13 == _T_973_0 ? _T_754_0_19 : _GEN_116;
  assign _GEN_118 = 5'h14 == _T_973_0 ? _T_754_0_20 : _GEN_117;
  assign _GEN_119 = 5'h15 == _T_973_0 ? _T_754_0_21 : _GEN_118;
  assign _GEN_120 = 5'h16 == _T_973_0 ? _T_754_0_22 : _GEN_119;
  assign _GEN_121 = 5'h17 == _T_973_0 ? _T_754_0_23 : _GEN_120;
  assign _GEN_122 = 5'h18 == _T_973_0 ? _T_754_0_24 : _GEN_121;
  assign _GEN_123 = 5'h19 == _T_973_0 ? _T_754_0_25 : _GEN_122;
  assign _GEN_124 = 5'h1a == _T_973_0 ? _T_754_0_26 : _GEN_123;
  assign _GEN_125 = 5'h1b == _T_973_0 ? _T_754_0_27 : _GEN_124;
  assign _GEN_126 = 5'h1c == _T_973_0 ? _T_754_0_28 : _GEN_125;
  assign _GEN_127 = 5'h1d == _T_973_0 ? _T_754_0_29 : _GEN_126;
  assign _GEN_128 = 5'h1e == _T_973_0 ? _T_754_0_30 : _GEN_127;
  assign _GEN_129 = 5'h1f == _T_973_0 ? _T_754_0_31 : _GEN_128;
  assign _T_4545 = _T_389 - 1'h1;
  assign _T_4546 = $unsigned(_T_4545);
  assign _T_4547 = _T_4546[0:0];
  assign _T_4548 = _T_4518 ? 1'h0 : _T_4547;
  assign _T_4550 = 1'h0 < _T_1007;
  assign _T_4551 = _T_4550 ? _T_389 : _T_4548;
  assign _T_4553 = _T_4551 == 1'h0;
  assign _T_4555 = _T_4553 ? _T_994_0 : 1'h0;
  assign _T_4934 = _T_4558 == 1'h0;
  assign _T_4936 = _T_4934 == 1'h0;
  assign _T_4938 = _T_4558 + 1'h1;
  assign _T_4939 = _T_4938[0:0];
  assign _GEN_130 = _T_4936 ? _T_4939 : _T_4558;
  assign _T_4946 = _T_4934 & _T_446_0;
  assign _T_4952 = _T_4572_0 == 1'h0;
  assign _T_4953 = _T_4946 & _T_4952;
  assign _T_4955 = io_axi_inputMemAddrValids_1 & io_axi_inputMemAddrReadys_1;
  assign _T_4960 = _T_4934 & _T_452_0;
  assign _T_4967 = _T_4960 & _T_4952;
  assign _T_4968 = _T_4955 | _T_4967;
  assign _GEN_131 = io_axi_inputMemAddrValids_1 ? 1'h1 : _T_4593_0;
  assign _T_4980 = _T_4924 == 1'h0;
  assign _T_4991 = _T_4924 + 1'h1;
  assign _T_4992 = _T_4991[0:0];
  assign _GEN_133 = _T_4980 ? 1'h0 : _GEN_130;
  assign _GEN_134 = _T_4980 ? 1'h0 : _T_4992;
  assign _GEN_135 = _T_4968 ? 1'h1 : _T_4572_0;
  assign _GEN_136 = _T_4968 ? _GEN_131 : _T_4593_0;
  assign _GEN_138 = _T_4968 ? _GEN_133 : _GEN_130;
  assign _GEN_139 = _T_4968 ? _GEN_134 : _T_4924;
  assign _T_4994 = _T_4893_0 == 5'h1f;
  assign _T_5000 = _T_4893_0 + 5'h1;
  assign _T_5001 = _T_5000[4:0];
  assign _GEN_140 = _T_4994 ? 1'h0 : _GEN_135;
  assign _GEN_141 = _T_4994 ? 1'h0 : _GEN_136;
  assign _GEN_142 = _T_4994 ? 1'h0 : _T_4914_0;
  assign _GEN_143 = _T_4994 ? 5'h0 : _T_5001;
  assign _GEN_144 = _T_4914_0 ? _GEN_140 : _GEN_135;
  assign _GEN_145 = _T_4914_0 ? _GEN_141 : _GEN_136;
  assign _GEN_146 = _T_4914_0 ? _GEN_142 : _T_4914_0;
  assign _GEN_147 = _T_4914_0 ? _GEN_143 : _T_4893_0;
  assign _T_5002 = io_axi_inputMemBlockReadys_1 & io_axi_inputMemBlockValids_1;
  assign _T_5007 = _T_4930 + 1'h1;
  assign _T_5008 = _T_5007[0:0];
  assign _T_5009 = _T_4930 ? 1'h0 : _T_5008;
  assign _T_5011 = 1'h0 == _T_4930;
  assign _T_5115 = io_axi_inputMemBlocks_1[31:0];
  assign _GEN_148 = _T_5011 ? _T_5115 : _T_4674_0_0;
  assign _T_5221 = io_axi_inputMemBlocks_1[63:32];
  assign _GEN_149 = _T_5011 ? _T_5221 : _T_4674_0_1;
  assign _T_5327 = io_axi_inputMemBlocks_1[95:64];
  assign _GEN_150 = _T_5011 ? _T_5327 : _T_4674_0_2;
  assign _T_5433 = io_axi_inputMemBlocks_1[127:96];
  assign _GEN_151 = _T_5011 ? _T_5433 : _T_4674_0_3;
  assign _T_5539 = io_axi_inputMemBlocks_1[159:128];
  assign _GEN_152 = _T_5011 ? _T_5539 : _T_4674_0_4;
  assign _T_5645 = io_axi_inputMemBlocks_1[191:160];
  assign _GEN_153 = _T_5011 ? _T_5645 : _T_4674_0_5;
  assign _T_5751 = io_axi_inputMemBlocks_1[223:192];
  assign _GEN_154 = _T_5011 ? _T_5751 : _T_4674_0_6;
  assign _T_5857 = io_axi_inputMemBlocks_1[255:224];
  assign _GEN_155 = _T_5011 ? _T_5857 : _T_4674_0_7;
  assign _T_5963 = io_axi_inputMemBlocks_1[287:256];
  assign _GEN_156 = _T_5011 ? _T_5963 : _T_4674_0_8;
  assign _T_6069 = io_axi_inputMemBlocks_1[319:288];
  assign _GEN_157 = _T_5011 ? _T_6069 : _T_4674_0_9;
  assign _T_6175 = io_axi_inputMemBlocks_1[351:320];
  assign _GEN_158 = _T_5011 ? _T_6175 : _T_4674_0_10;
  assign _T_6281 = io_axi_inputMemBlocks_1[383:352];
  assign _GEN_159 = _T_5011 ? _T_6281 : _T_4674_0_11;
  assign _T_6387 = io_axi_inputMemBlocks_1[415:384];
  assign _GEN_160 = _T_5011 ? _T_6387 : _T_4674_0_12;
  assign _T_6493 = io_axi_inputMemBlocks_1[447:416];
  assign _GEN_161 = _T_5011 ? _T_6493 : _T_4674_0_13;
  assign _T_6599 = io_axi_inputMemBlocks_1[479:448];
  assign _GEN_162 = _T_5011 ? _T_6599 : _T_4674_0_14;
  assign _T_6705 = io_axi_inputMemBlocks_1[511:480];
  assign _GEN_163 = _T_5011 ? _T_6705 : _T_4674_0_15;
  assign _GEN_164 = _T_4930 ? _T_5115 : _T_4674_0_16;
  assign _GEN_165 = _T_4930 ? _T_5221 : _T_4674_0_17;
  assign _GEN_166 = _T_4930 ? _T_5327 : _T_4674_0_18;
  assign _GEN_167 = _T_4930 ? _T_5433 : _T_4674_0_19;
  assign _GEN_168 = _T_4930 ? _T_5539 : _T_4674_0_20;
  assign _GEN_169 = _T_4930 ? _T_5645 : _T_4674_0_21;
  assign _GEN_170 = _T_4930 ? _T_5751 : _T_4674_0_22;
  assign _GEN_171 = _T_4930 ? _T_5857 : _T_4674_0_23;
  assign _GEN_172 = _T_4930 ? _T_5963 : _T_4674_0_24;
  assign _GEN_173 = _T_4930 ? _T_6069 : _T_4674_0_25;
  assign _GEN_174 = _T_4930 ? _T_6175 : _T_4674_0_26;
  assign _GEN_175 = _T_4930 ? _T_6281 : _T_4674_0_27;
  assign _GEN_176 = _T_4930 ? _T_6387 : _T_4674_0_28;
  assign _GEN_177 = _T_4930 ? _T_6493 : _T_4674_0_29;
  assign _GEN_178 = _T_4930 ? _T_6599 : _T_4674_0_30;
  assign _GEN_179 = _T_4930 ? _T_6705 : _T_4674_0_31;
  assign _GEN_180 = _T_5002 ? _T_5009 : _T_4930;
  assign _GEN_181 = _T_5002 ? _GEN_148 : _T_4674_0_0;
  assign _GEN_182 = _T_5002 ? _GEN_149 : _T_4674_0_1;
  assign _GEN_183 = _T_5002 ? _GEN_150 : _T_4674_0_2;
  assign _GEN_184 = _T_5002 ? _GEN_151 : _T_4674_0_3;
  assign _GEN_185 = _T_5002 ? _GEN_152 : _T_4674_0_4;
  assign _GEN_186 = _T_5002 ? _GEN_153 : _T_4674_0_5;
  assign _GEN_187 = _T_5002 ? _GEN_154 : _T_4674_0_6;
  assign _GEN_188 = _T_5002 ? _GEN_155 : _T_4674_0_7;
  assign _GEN_189 = _T_5002 ? _GEN_156 : _T_4674_0_8;
  assign _GEN_190 = _T_5002 ? _GEN_157 : _T_4674_0_9;
  assign _GEN_191 = _T_5002 ? _GEN_158 : _T_4674_0_10;
  assign _GEN_192 = _T_5002 ? _GEN_159 : _T_4674_0_11;
  assign _GEN_193 = _T_5002 ? _GEN_160 : _T_4674_0_12;
  assign _GEN_194 = _T_5002 ? _GEN_161 : _T_4674_0_13;
  assign _GEN_195 = _T_5002 ? _GEN_162 : _T_4674_0_14;
  assign _GEN_196 = _T_5002 ? _GEN_163 : _T_4674_0_15;
  assign _GEN_197 = _T_5002 ? _GEN_164 : _T_4674_0_16;
  assign _GEN_198 = _T_5002 ? _GEN_165 : _T_4674_0_17;
  assign _GEN_199 = _T_5002 ? _GEN_166 : _T_4674_0_18;
  assign _GEN_200 = _T_5002 ? _GEN_167 : _T_4674_0_19;
  assign _GEN_201 = _T_5002 ? _GEN_168 : _T_4674_0_20;
  assign _GEN_202 = _T_5002 ? _GEN_169 : _T_4674_0_21;
  assign _GEN_203 = _T_5002 ? _GEN_170 : _T_4674_0_22;
  assign _GEN_204 = _T_5002 ? _GEN_171 : _T_4674_0_23;
  assign _GEN_205 = _T_5002 ? _GEN_172 : _T_4674_0_24;
  assign _GEN_206 = _T_5002 ? _GEN_173 : _T_4674_0_25;
  assign _GEN_207 = _T_5002 ? _GEN_174 : _T_4674_0_26;
  assign _GEN_208 = _T_5002 ? _GEN_175 : _T_4674_0_27;
  assign _GEN_209 = _T_5002 ? _GEN_176 : _T_4674_0_28;
  assign _GEN_210 = _T_5002 ? _GEN_177 : _T_4674_0_29;
  assign _GEN_211 = _T_5002 ? _GEN_178 : _T_4674_0_30;
  assign _GEN_212 = _T_5002 ? _GEN_179 : _T_4674_0_31;
  assign _T_8402 = io_axi_inputMemBlockValids_1 & io_axi_inputMemBlockReadys_1;
  assign _T_8405 = _T_8402 & _T_4930;
  assign _T_8415 = _T_4593_0 == 1'h0;
  assign _T_8416 = _T_4572_0 & _T_8415;
  assign _T_8422 = _T_4914_0 == 1'h0;
  assign _T_8423 = _T_8416 & _T_8422;
  assign _T_8424 = _T_8405 | _T_8423;
  assign _GEN_213 = io_axi_inputMemBlockReadys_1 ? 1'h1 : _GEN_146;
  assign _GEN_214 = io_axi_inputMemBlockReadys_1 ? _GEN_144 : 1'h0;
  assign _T_8436 = _T_4927 == 1'h0;
  assign _T_8438 = _T_395 == 1'h0;
  assign _T_8441 = _T_395 + 1'h1;
  assign _T_8442 = _T_8441[0:0];
  assign _T_8443 = _T_8438 ? 1'h0 : _T_8442;
  assign _T_8446 = _T_4927 + 1'h1;
  assign _T_8447 = _T_8446[0:0];
  assign _GEN_215 = _T_8436 ? _T_8443 : _T_395;
  assign _GEN_216 = _T_8436 ? 1'h0 : _T_8447;
  assign _GEN_217 = _T_8424 ? _GEN_213 : _GEN_146;
  assign _GEN_218 = _T_8424 ? _GEN_214 : _GEN_144;
  assign _GEN_219 = _T_8424 ? _GEN_215 : _T_395;
  assign _GEN_220 = _T_8424 ? _GEN_216 : _T_4927;
  assign _T_8458 = _T_4593_0 & _T_8422;
  assign _GEN_221 = 5'h1 == _T_4893_0 ? _T_4674_0_1 : _T_4674_0_0;
  assign _GEN_222 = 5'h2 == _T_4893_0 ? _T_4674_0_2 : _GEN_221;
  assign _GEN_223 = 5'h3 == _T_4893_0 ? _T_4674_0_3 : _GEN_222;
  assign _GEN_224 = 5'h4 == _T_4893_0 ? _T_4674_0_4 : _GEN_223;
  assign _GEN_225 = 5'h5 == _T_4893_0 ? _T_4674_0_5 : _GEN_224;
  assign _GEN_226 = 5'h6 == _T_4893_0 ? _T_4674_0_6 : _GEN_225;
  assign _GEN_227 = 5'h7 == _T_4893_0 ? _T_4674_0_7 : _GEN_226;
  assign _GEN_228 = 5'h8 == _T_4893_0 ? _T_4674_0_8 : _GEN_227;
  assign _GEN_229 = 5'h9 == _T_4893_0 ? _T_4674_0_9 : _GEN_228;
  assign _GEN_230 = 5'ha == _T_4893_0 ? _T_4674_0_10 : _GEN_229;
  assign _GEN_231 = 5'hb == _T_4893_0 ? _T_4674_0_11 : _GEN_230;
  assign _GEN_232 = 5'hc == _T_4893_0 ? _T_4674_0_12 : _GEN_231;
  assign _GEN_233 = 5'hd == _T_4893_0 ? _T_4674_0_13 : _GEN_232;
  assign _GEN_234 = 5'he == _T_4893_0 ? _T_4674_0_14 : _GEN_233;
  assign _GEN_235 = 5'hf == _T_4893_0 ? _T_4674_0_15 : _GEN_234;
  assign _GEN_236 = 5'h10 == _T_4893_0 ? _T_4674_0_16 : _GEN_235;
  assign _GEN_237 = 5'h11 == _T_4893_0 ? _T_4674_0_17 : _GEN_236;
  assign _GEN_238 = 5'h12 == _T_4893_0 ? _T_4674_0_18 : _GEN_237;
  assign _GEN_239 = 5'h13 == _T_4893_0 ? _T_4674_0_19 : _GEN_238;
  assign _GEN_240 = 5'h14 == _T_4893_0 ? _T_4674_0_20 : _GEN_239;
  assign _GEN_241 = 5'h15 == _T_4893_0 ? _T_4674_0_21 : _GEN_240;
  assign _GEN_242 = 5'h16 == _T_4893_0 ? _T_4674_0_22 : _GEN_241;
  assign _GEN_243 = 5'h17 == _T_4893_0 ? _T_4674_0_23 : _GEN_242;
  assign _GEN_244 = 5'h18 == _T_4893_0 ? _T_4674_0_24 : _GEN_243;
  assign _GEN_245 = 5'h19 == _T_4893_0 ? _T_4674_0_25 : _GEN_244;
  assign _GEN_246 = 5'h1a == _T_4893_0 ? _T_4674_0_26 : _GEN_245;
  assign _GEN_247 = 5'h1b == _T_4893_0 ? _T_4674_0_27 : _GEN_246;
  assign _GEN_248 = 5'h1c == _T_4893_0 ? _T_4674_0_28 : _GEN_247;
  assign _GEN_249 = 5'h1d == _T_4893_0 ? _T_4674_0_29 : _GEN_248;
  assign _GEN_250 = 5'h1e == _T_4893_0 ? _T_4674_0_30 : _GEN_249;
  assign _GEN_251 = 5'h1f == _T_4893_0 ? _T_4674_0_31 : _GEN_250;
  assign _T_8465 = _T_395 - 1'h1;
  assign _T_8466 = $unsigned(_T_8465);
  assign _T_8467 = _T_8466[0:0];
  assign _T_8468 = _T_8438 ? 1'h0 : _T_8467;
  assign _T_8470 = 1'h0 < _T_4927;
  assign _T_8471 = _T_8470 ? _T_395 : _T_8468;
  assign _T_8473 = _T_8471 == 1'h0;
  assign _T_8475 = _T_8473 ? _T_4914_0 : 1'h0;
  assign _T_8854 = _T_8478 == 1'h0;
  assign _T_8856 = _T_8854 == 1'h0;
  assign _T_8858 = _T_8478 + 1'h1;
  assign _T_8859 = _T_8858[0:0];
  assign _GEN_252 = _T_8856 ? _T_8859 : _T_8478;
  assign _T_8866 = _T_8854 & _T_464_0;
  assign _T_8872 = _T_8492_0 == 1'h0;
  assign _T_8873 = _T_8866 & _T_8872;
  assign _T_8875 = io_axi_inputMemAddrValids_2 & io_axi_inputMemAddrReadys_2;
  assign _T_8880 = _T_8854 & _T_470_0;
  assign _T_8887 = _T_8880 & _T_8872;
  assign _T_8888 = _T_8875 | _T_8887;
  assign _GEN_253 = io_axi_inputMemAddrValids_2 ? 1'h1 : _T_8513_0;
  assign _T_8900 = _T_8844 == 1'h0;
  assign _T_8911 = _T_8844 + 1'h1;
  assign _T_8912 = _T_8911[0:0];
  assign _GEN_255 = _T_8900 ? 1'h0 : _GEN_252;
  assign _GEN_256 = _T_8900 ? 1'h0 : _T_8912;
  assign _GEN_257 = _T_8888 ? 1'h1 : _T_8492_0;
  assign _GEN_258 = _T_8888 ? _GEN_253 : _T_8513_0;
  assign _GEN_260 = _T_8888 ? _GEN_255 : _GEN_252;
  assign _GEN_261 = _T_8888 ? _GEN_256 : _T_8844;
  assign _T_8914 = _T_8813_0 == 5'h1f;
  assign _T_8920 = _T_8813_0 + 5'h1;
  assign _T_8921 = _T_8920[4:0];
  assign _GEN_262 = _T_8914 ? 1'h0 : _GEN_257;
  assign _GEN_263 = _T_8914 ? 1'h0 : _GEN_258;
  assign _GEN_264 = _T_8914 ? 1'h0 : _T_8834_0;
  assign _GEN_265 = _T_8914 ? 5'h0 : _T_8921;
  assign _GEN_266 = _T_8834_0 ? _GEN_262 : _GEN_257;
  assign _GEN_267 = _T_8834_0 ? _GEN_263 : _GEN_258;
  assign _GEN_268 = _T_8834_0 ? _GEN_264 : _T_8834_0;
  assign _GEN_269 = _T_8834_0 ? _GEN_265 : _T_8813_0;
  assign _T_8922 = io_axi_inputMemBlockReadys_2 & io_axi_inputMemBlockValids_2;
  assign _T_8927 = _T_8850 + 1'h1;
  assign _T_8928 = _T_8927[0:0];
  assign _T_8929 = _T_8850 ? 1'h0 : _T_8928;
  assign _T_8931 = 1'h0 == _T_8850;
  assign _T_9035 = io_axi_inputMemBlocks_2[31:0];
  assign _GEN_270 = _T_8931 ? _T_9035 : _T_8594_0_0;
  assign _T_9141 = io_axi_inputMemBlocks_2[63:32];
  assign _GEN_271 = _T_8931 ? _T_9141 : _T_8594_0_1;
  assign _T_9247 = io_axi_inputMemBlocks_2[95:64];
  assign _GEN_272 = _T_8931 ? _T_9247 : _T_8594_0_2;
  assign _T_9353 = io_axi_inputMemBlocks_2[127:96];
  assign _GEN_273 = _T_8931 ? _T_9353 : _T_8594_0_3;
  assign _T_9459 = io_axi_inputMemBlocks_2[159:128];
  assign _GEN_274 = _T_8931 ? _T_9459 : _T_8594_0_4;
  assign _T_9565 = io_axi_inputMemBlocks_2[191:160];
  assign _GEN_275 = _T_8931 ? _T_9565 : _T_8594_0_5;
  assign _T_9671 = io_axi_inputMemBlocks_2[223:192];
  assign _GEN_276 = _T_8931 ? _T_9671 : _T_8594_0_6;
  assign _T_9777 = io_axi_inputMemBlocks_2[255:224];
  assign _GEN_277 = _T_8931 ? _T_9777 : _T_8594_0_7;
  assign _T_9883 = io_axi_inputMemBlocks_2[287:256];
  assign _GEN_278 = _T_8931 ? _T_9883 : _T_8594_0_8;
  assign _T_9989 = io_axi_inputMemBlocks_2[319:288];
  assign _GEN_279 = _T_8931 ? _T_9989 : _T_8594_0_9;
  assign _T_10095 = io_axi_inputMemBlocks_2[351:320];
  assign _GEN_280 = _T_8931 ? _T_10095 : _T_8594_0_10;
  assign _T_10201 = io_axi_inputMemBlocks_2[383:352];
  assign _GEN_281 = _T_8931 ? _T_10201 : _T_8594_0_11;
  assign _T_10307 = io_axi_inputMemBlocks_2[415:384];
  assign _GEN_282 = _T_8931 ? _T_10307 : _T_8594_0_12;
  assign _T_10413 = io_axi_inputMemBlocks_2[447:416];
  assign _GEN_283 = _T_8931 ? _T_10413 : _T_8594_0_13;
  assign _T_10519 = io_axi_inputMemBlocks_2[479:448];
  assign _GEN_284 = _T_8931 ? _T_10519 : _T_8594_0_14;
  assign _T_10625 = io_axi_inputMemBlocks_2[511:480];
  assign _GEN_285 = _T_8931 ? _T_10625 : _T_8594_0_15;
  assign _GEN_286 = _T_8850 ? _T_9035 : _T_8594_0_16;
  assign _GEN_287 = _T_8850 ? _T_9141 : _T_8594_0_17;
  assign _GEN_288 = _T_8850 ? _T_9247 : _T_8594_0_18;
  assign _GEN_289 = _T_8850 ? _T_9353 : _T_8594_0_19;
  assign _GEN_290 = _T_8850 ? _T_9459 : _T_8594_0_20;
  assign _GEN_291 = _T_8850 ? _T_9565 : _T_8594_0_21;
  assign _GEN_292 = _T_8850 ? _T_9671 : _T_8594_0_22;
  assign _GEN_293 = _T_8850 ? _T_9777 : _T_8594_0_23;
  assign _GEN_294 = _T_8850 ? _T_9883 : _T_8594_0_24;
  assign _GEN_295 = _T_8850 ? _T_9989 : _T_8594_0_25;
  assign _GEN_296 = _T_8850 ? _T_10095 : _T_8594_0_26;
  assign _GEN_297 = _T_8850 ? _T_10201 : _T_8594_0_27;
  assign _GEN_298 = _T_8850 ? _T_10307 : _T_8594_0_28;
  assign _GEN_299 = _T_8850 ? _T_10413 : _T_8594_0_29;
  assign _GEN_300 = _T_8850 ? _T_10519 : _T_8594_0_30;
  assign _GEN_301 = _T_8850 ? _T_10625 : _T_8594_0_31;
  assign _GEN_302 = _T_8922 ? _T_8929 : _T_8850;
  assign _GEN_303 = _T_8922 ? _GEN_270 : _T_8594_0_0;
  assign _GEN_304 = _T_8922 ? _GEN_271 : _T_8594_0_1;
  assign _GEN_305 = _T_8922 ? _GEN_272 : _T_8594_0_2;
  assign _GEN_306 = _T_8922 ? _GEN_273 : _T_8594_0_3;
  assign _GEN_307 = _T_8922 ? _GEN_274 : _T_8594_0_4;
  assign _GEN_308 = _T_8922 ? _GEN_275 : _T_8594_0_5;
  assign _GEN_309 = _T_8922 ? _GEN_276 : _T_8594_0_6;
  assign _GEN_310 = _T_8922 ? _GEN_277 : _T_8594_0_7;
  assign _GEN_311 = _T_8922 ? _GEN_278 : _T_8594_0_8;
  assign _GEN_312 = _T_8922 ? _GEN_279 : _T_8594_0_9;
  assign _GEN_313 = _T_8922 ? _GEN_280 : _T_8594_0_10;
  assign _GEN_314 = _T_8922 ? _GEN_281 : _T_8594_0_11;
  assign _GEN_315 = _T_8922 ? _GEN_282 : _T_8594_0_12;
  assign _GEN_316 = _T_8922 ? _GEN_283 : _T_8594_0_13;
  assign _GEN_317 = _T_8922 ? _GEN_284 : _T_8594_0_14;
  assign _GEN_318 = _T_8922 ? _GEN_285 : _T_8594_0_15;
  assign _GEN_319 = _T_8922 ? _GEN_286 : _T_8594_0_16;
  assign _GEN_320 = _T_8922 ? _GEN_287 : _T_8594_0_17;
  assign _GEN_321 = _T_8922 ? _GEN_288 : _T_8594_0_18;
  assign _GEN_322 = _T_8922 ? _GEN_289 : _T_8594_0_19;
  assign _GEN_323 = _T_8922 ? _GEN_290 : _T_8594_0_20;
  assign _GEN_324 = _T_8922 ? _GEN_291 : _T_8594_0_21;
  assign _GEN_325 = _T_8922 ? _GEN_292 : _T_8594_0_22;
  assign _GEN_326 = _T_8922 ? _GEN_293 : _T_8594_0_23;
  assign _GEN_327 = _T_8922 ? _GEN_294 : _T_8594_0_24;
  assign _GEN_328 = _T_8922 ? _GEN_295 : _T_8594_0_25;
  assign _GEN_329 = _T_8922 ? _GEN_296 : _T_8594_0_26;
  assign _GEN_330 = _T_8922 ? _GEN_297 : _T_8594_0_27;
  assign _GEN_331 = _T_8922 ? _GEN_298 : _T_8594_0_28;
  assign _GEN_332 = _T_8922 ? _GEN_299 : _T_8594_0_29;
  assign _GEN_333 = _T_8922 ? _GEN_300 : _T_8594_0_30;
  assign _GEN_334 = _T_8922 ? _GEN_301 : _T_8594_0_31;
  assign _T_12322 = io_axi_inputMemBlockValids_2 & io_axi_inputMemBlockReadys_2;
  assign _T_12325 = _T_12322 & _T_8850;
  assign _T_12335 = _T_8513_0 == 1'h0;
  assign _T_12336 = _T_8492_0 & _T_12335;
  assign _T_12342 = _T_8834_0 == 1'h0;
  assign _T_12343 = _T_12336 & _T_12342;
  assign _T_12344 = _T_12325 | _T_12343;
  assign _GEN_335 = io_axi_inputMemBlockReadys_2 ? 1'h1 : _GEN_268;
  assign _GEN_336 = io_axi_inputMemBlockReadys_2 ? _GEN_266 : 1'h0;
  assign _T_12356 = _T_8847 == 1'h0;
  assign _T_12358 = _T_401 == 1'h0;
  assign _T_12361 = _T_401 + 1'h1;
  assign _T_12362 = _T_12361[0:0];
  assign _T_12363 = _T_12358 ? 1'h0 : _T_12362;
  assign _T_12366 = _T_8847 + 1'h1;
  assign _T_12367 = _T_12366[0:0];
  assign _GEN_337 = _T_12356 ? _T_12363 : _T_401;
  assign _GEN_338 = _T_12356 ? 1'h0 : _T_12367;
  assign _GEN_339 = _T_12344 ? _GEN_335 : _GEN_268;
  assign _GEN_340 = _T_12344 ? _GEN_336 : _GEN_266;
  assign _GEN_341 = _T_12344 ? _GEN_337 : _T_401;
  assign _GEN_342 = _T_12344 ? _GEN_338 : _T_8847;
  assign _T_12378 = _T_8513_0 & _T_12342;
  assign _GEN_343 = 5'h1 == _T_8813_0 ? _T_8594_0_1 : _T_8594_0_0;
  assign _GEN_344 = 5'h2 == _T_8813_0 ? _T_8594_0_2 : _GEN_343;
  assign _GEN_345 = 5'h3 == _T_8813_0 ? _T_8594_0_3 : _GEN_344;
  assign _GEN_346 = 5'h4 == _T_8813_0 ? _T_8594_0_4 : _GEN_345;
  assign _GEN_347 = 5'h5 == _T_8813_0 ? _T_8594_0_5 : _GEN_346;
  assign _GEN_348 = 5'h6 == _T_8813_0 ? _T_8594_0_6 : _GEN_347;
  assign _GEN_349 = 5'h7 == _T_8813_0 ? _T_8594_0_7 : _GEN_348;
  assign _GEN_350 = 5'h8 == _T_8813_0 ? _T_8594_0_8 : _GEN_349;
  assign _GEN_351 = 5'h9 == _T_8813_0 ? _T_8594_0_9 : _GEN_350;
  assign _GEN_352 = 5'ha == _T_8813_0 ? _T_8594_0_10 : _GEN_351;
  assign _GEN_353 = 5'hb == _T_8813_0 ? _T_8594_0_11 : _GEN_352;
  assign _GEN_354 = 5'hc == _T_8813_0 ? _T_8594_0_12 : _GEN_353;
  assign _GEN_355 = 5'hd == _T_8813_0 ? _T_8594_0_13 : _GEN_354;
  assign _GEN_356 = 5'he == _T_8813_0 ? _T_8594_0_14 : _GEN_355;
  assign _GEN_357 = 5'hf == _T_8813_0 ? _T_8594_0_15 : _GEN_356;
  assign _GEN_358 = 5'h10 == _T_8813_0 ? _T_8594_0_16 : _GEN_357;
  assign _GEN_359 = 5'h11 == _T_8813_0 ? _T_8594_0_17 : _GEN_358;
  assign _GEN_360 = 5'h12 == _T_8813_0 ? _T_8594_0_18 : _GEN_359;
  assign _GEN_361 = 5'h13 == _T_8813_0 ? _T_8594_0_19 : _GEN_360;
  assign _GEN_362 = 5'h14 == _T_8813_0 ? _T_8594_0_20 : _GEN_361;
  assign _GEN_363 = 5'h15 == _T_8813_0 ? _T_8594_0_21 : _GEN_362;
  assign _GEN_364 = 5'h16 == _T_8813_0 ? _T_8594_0_22 : _GEN_363;
  assign _GEN_365 = 5'h17 == _T_8813_0 ? _T_8594_0_23 : _GEN_364;
  assign _GEN_366 = 5'h18 == _T_8813_0 ? _T_8594_0_24 : _GEN_365;
  assign _GEN_367 = 5'h19 == _T_8813_0 ? _T_8594_0_25 : _GEN_366;
  assign _GEN_368 = 5'h1a == _T_8813_0 ? _T_8594_0_26 : _GEN_367;
  assign _GEN_369 = 5'h1b == _T_8813_0 ? _T_8594_0_27 : _GEN_368;
  assign _GEN_370 = 5'h1c == _T_8813_0 ? _T_8594_0_28 : _GEN_369;
  assign _GEN_371 = 5'h1d == _T_8813_0 ? _T_8594_0_29 : _GEN_370;
  assign _GEN_372 = 5'h1e == _T_8813_0 ? _T_8594_0_30 : _GEN_371;
  assign _GEN_373 = 5'h1f == _T_8813_0 ? _T_8594_0_31 : _GEN_372;
  assign _T_12385 = _T_401 - 1'h1;
  assign _T_12386 = $unsigned(_T_12385);
  assign _T_12387 = _T_12386[0:0];
  assign _T_12388 = _T_12358 ? 1'h0 : _T_12387;
  assign _T_12390 = 1'h0 < _T_8847;
  assign _T_12391 = _T_12390 ? _T_401 : _T_12388;
  assign _T_12393 = _T_12391 == 1'h0;
  assign _T_12395 = _T_12393 ? _T_8834_0 : 1'h0;
  assign _T_12774 = _T_12398 == 1'h0;
  assign _T_12776 = _T_12774 == 1'h0;
  assign _T_12778 = _T_12398 + 1'h1;
  assign _T_12779 = _T_12778[0:0];
  assign _GEN_374 = _T_12776 ? _T_12779 : _T_12398;
  assign _T_12786 = _T_12774 & _T_482_0;
  assign _T_12792 = _T_12412_0 == 1'h0;
  assign _T_12793 = _T_12786 & _T_12792;
  assign _T_12795 = io_axi_inputMemAddrValids_3 & io_axi_inputMemAddrReadys_3;
  assign _T_12800 = _T_12774 & _T_488_0;
  assign _T_12807 = _T_12800 & _T_12792;
  assign _T_12808 = _T_12795 | _T_12807;
  assign _GEN_375 = io_axi_inputMemAddrValids_3 ? 1'h1 : _T_12433_0;
  assign _T_12820 = _T_12764 == 1'h0;
  assign _T_12831 = _T_12764 + 1'h1;
  assign _T_12832 = _T_12831[0:0];
  assign _GEN_377 = _T_12820 ? 1'h0 : _GEN_374;
  assign _GEN_378 = _T_12820 ? 1'h0 : _T_12832;
  assign _GEN_379 = _T_12808 ? 1'h1 : _T_12412_0;
  assign _GEN_380 = _T_12808 ? _GEN_375 : _T_12433_0;
  assign _GEN_382 = _T_12808 ? _GEN_377 : _GEN_374;
  assign _GEN_383 = _T_12808 ? _GEN_378 : _T_12764;
  assign _T_12834 = _T_12733_0 == 5'h1f;
  assign _T_12840 = _T_12733_0 + 5'h1;
  assign _T_12841 = _T_12840[4:0];
  assign _GEN_384 = _T_12834 ? 1'h0 : _GEN_379;
  assign _GEN_385 = _T_12834 ? 1'h0 : _GEN_380;
  assign _GEN_386 = _T_12834 ? 1'h0 : _T_12754_0;
  assign _GEN_387 = _T_12834 ? 5'h0 : _T_12841;
  assign _GEN_388 = _T_12754_0 ? _GEN_384 : _GEN_379;
  assign _GEN_389 = _T_12754_0 ? _GEN_385 : _GEN_380;
  assign _GEN_390 = _T_12754_0 ? _GEN_386 : _T_12754_0;
  assign _GEN_391 = _T_12754_0 ? _GEN_387 : _T_12733_0;
  assign _T_12842 = io_axi_inputMemBlockReadys_3 & io_axi_inputMemBlockValids_3;
  assign _T_12847 = _T_12770 + 1'h1;
  assign _T_12848 = _T_12847[0:0];
  assign _T_12849 = _T_12770 ? 1'h0 : _T_12848;
  assign _T_12851 = 1'h0 == _T_12770;
  assign _T_12955 = io_axi_inputMemBlocks_3[31:0];
  assign _GEN_392 = _T_12851 ? _T_12955 : _T_12514_0_0;
  assign _T_13061 = io_axi_inputMemBlocks_3[63:32];
  assign _GEN_393 = _T_12851 ? _T_13061 : _T_12514_0_1;
  assign _T_13167 = io_axi_inputMemBlocks_3[95:64];
  assign _GEN_394 = _T_12851 ? _T_13167 : _T_12514_0_2;
  assign _T_13273 = io_axi_inputMemBlocks_3[127:96];
  assign _GEN_395 = _T_12851 ? _T_13273 : _T_12514_0_3;
  assign _T_13379 = io_axi_inputMemBlocks_3[159:128];
  assign _GEN_396 = _T_12851 ? _T_13379 : _T_12514_0_4;
  assign _T_13485 = io_axi_inputMemBlocks_3[191:160];
  assign _GEN_397 = _T_12851 ? _T_13485 : _T_12514_0_5;
  assign _T_13591 = io_axi_inputMemBlocks_3[223:192];
  assign _GEN_398 = _T_12851 ? _T_13591 : _T_12514_0_6;
  assign _T_13697 = io_axi_inputMemBlocks_3[255:224];
  assign _GEN_399 = _T_12851 ? _T_13697 : _T_12514_0_7;
  assign _T_13803 = io_axi_inputMemBlocks_3[287:256];
  assign _GEN_400 = _T_12851 ? _T_13803 : _T_12514_0_8;
  assign _T_13909 = io_axi_inputMemBlocks_3[319:288];
  assign _GEN_401 = _T_12851 ? _T_13909 : _T_12514_0_9;
  assign _T_14015 = io_axi_inputMemBlocks_3[351:320];
  assign _GEN_402 = _T_12851 ? _T_14015 : _T_12514_0_10;
  assign _T_14121 = io_axi_inputMemBlocks_3[383:352];
  assign _GEN_403 = _T_12851 ? _T_14121 : _T_12514_0_11;
  assign _T_14227 = io_axi_inputMemBlocks_3[415:384];
  assign _GEN_404 = _T_12851 ? _T_14227 : _T_12514_0_12;
  assign _T_14333 = io_axi_inputMemBlocks_3[447:416];
  assign _GEN_405 = _T_12851 ? _T_14333 : _T_12514_0_13;
  assign _T_14439 = io_axi_inputMemBlocks_3[479:448];
  assign _GEN_406 = _T_12851 ? _T_14439 : _T_12514_0_14;
  assign _T_14545 = io_axi_inputMemBlocks_3[511:480];
  assign _GEN_407 = _T_12851 ? _T_14545 : _T_12514_0_15;
  assign _GEN_408 = _T_12770 ? _T_12955 : _T_12514_0_16;
  assign _GEN_409 = _T_12770 ? _T_13061 : _T_12514_0_17;
  assign _GEN_410 = _T_12770 ? _T_13167 : _T_12514_0_18;
  assign _GEN_411 = _T_12770 ? _T_13273 : _T_12514_0_19;
  assign _GEN_412 = _T_12770 ? _T_13379 : _T_12514_0_20;
  assign _GEN_413 = _T_12770 ? _T_13485 : _T_12514_0_21;
  assign _GEN_414 = _T_12770 ? _T_13591 : _T_12514_0_22;
  assign _GEN_415 = _T_12770 ? _T_13697 : _T_12514_0_23;
  assign _GEN_416 = _T_12770 ? _T_13803 : _T_12514_0_24;
  assign _GEN_417 = _T_12770 ? _T_13909 : _T_12514_0_25;
  assign _GEN_418 = _T_12770 ? _T_14015 : _T_12514_0_26;
  assign _GEN_419 = _T_12770 ? _T_14121 : _T_12514_0_27;
  assign _GEN_420 = _T_12770 ? _T_14227 : _T_12514_0_28;
  assign _GEN_421 = _T_12770 ? _T_14333 : _T_12514_0_29;
  assign _GEN_422 = _T_12770 ? _T_14439 : _T_12514_0_30;
  assign _GEN_423 = _T_12770 ? _T_14545 : _T_12514_0_31;
  assign _GEN_424 = _T_12842 ? _T_12849 : _T_12770;
  assign _GEN_425 = _T_12842 ? _GEN_392 : _T_12514_0_0;
  assign _GEN_426 = _T_12842 ? _GEN_393 : _T_12514_0_1;
  assign _GEN_427 = _T_12842 ? _GEN_394 : _T_12514_0_2;
  assign _GEN_428 = _T_12842 ? _GEN_395 : _T_12514_0_3;
  assign _GEN_429 = _T_12842 ? _GEN_396 : _T_12514_0_4;
  assign _GEN_430 = _T_12842 ? _GEN_397 : _T_12514_0_5;
  assign _GEN_431 = _T_12842 ? _GEN_398 : _T_12514_0_6;
  assign _GEN_432 = _T_12842 ? _GEN_399 : _T_12514_0_7;
  assign _GEN_433 = _T_12842 ? _GEN_400 : _T_12514_0_8;
  assign _GEN_434 = _T_12842 ? _GEN_401 : _T_12514_0_9;
  assign _GEN_435 = _T_12842 ? _GEN_402 : _T_12514_0_10;
  assign _GEN_436 = _T_12842 ? _GEN_403 : _T_12514_0_11;
  assign _GEN_437 = _T_12842 ? _GEN_404 : _T_12514_0_12;
  assign _GEN_438 = _T_12842 ? _GEN_405 : _T_12514_0_13;
  assign _GEN_439 = _T_12842 ? _GEN_406 : _T_12514_0_14;
  assign _GEN_440 = _T_12842 ? _GEN_407 : _T_12514_0_15;
  assign _GEN_441 = _T_12842 ? _GEN_408 : _T_12514_0_16;
  assign _GEN_442 = _T_12842 ? _GEN_409 : _T_12514_0_17;
  assign _GEN_443 = _T_12842 ? _GEN_410 : _T_12514_0_18;
  assign _GEN_444 = _T_12842 ? _GEN_411 : _T_12514_0_19;
  assign _GEN_445 = _T_12842 ? _GEN_412 : _T_12514_0_20;
  assign _GEN_446 = _T_12842 ? _GEN_413 : _T_12514_0_21;
  assign _GEN_447 = _T_12842 ? _GEN_414 : _T_12514_0_22;
  assign _GEN_448 = _T_12842 ? _GEN_415 : _T_12514_0_23;
  assign _GEN_449 = _T_12842 ? _GEN_416 : _T_12514_0_24;
  assign _GEN_450 = _T_12842 ? _GEN_417 : _T_12514_0_25;
  assign _GEN_451 = _T_12842 ? _GEN_418 : _T_12514_0_26;
  assign _GEN_452 = _T_12842 ? _GEN_419 : _T_12514_0_27;
  assign _GEN_453 = _T_12842 ? _GEN_420 : _T_12514_0_28;
  assign _GEN_454 = _T_12842 ? _GEN_421 : _T_12514_0_29;
  assign _GEN_455 = _T_12842 ? _GEN_422 : _T_12514_0_30;
  assign _GEN_456 = _T_12842 ? _GEN_423 : _T_12514_0_31;
  assign _T_16242 = io_axi_inputMemBlockValids_3 & io_axi_inputMemBlockReadys_3;
  assign _T_16245 = _T_16242 & _T_12770;
  assign _T_16255 = _T_12433_0 == 1'h0;
  assign _T_16256 = _T_12412_0 & _T_16255;
  assign _T_16262 = _T_12754_0 == 1'h0;
  assign _T_16263 = _T_16256 & _T_16262;
  assign _T_16264 = _T_16245 | _T_16263;
  assign _GEN_457 = io_axi_inputMemBlockReadys_3 ? 1'h1 : _GEN_390;
  assign _GEN_458 = io_axi_inputMemBlockReadys_3 ? _GEN_388 : 1'h0;
  assign _T_16276 = _T_12767 == 1'h0;
  assign _T_16278 = _T_407 == 1'h0;
  assign _T_16281 = _T_407 + 1'h1;
  assign _T_16282 = _T_16281[0:0];
  assign _T_16283 = _T_16278 ? 1'h0 : _T_16282;
  assign _T_16286 = _T_12767 + 1'h1;
  assign _T_16287 = _T_16286[0:0];
  assign _GEN_459 = _T_16276 ? _T_16283 : _T_407;
  assign _GEN_460 = _T_16276 ? 1'h0 : _T_16287;
  assign _GEN_461 = _T_16264 ? _GEN_457 : _GEN_390;
  assign _GEN_462 = _T_16264 ? _GEN_458 : _GEN_388;
  assign _GEN_463 = _T_16264 ? _GEN_459 : _T_407;
  assign _GEN_464 = _T_16264 ? _GEN_460 : _T_12767;
  assign _T_16298 = _T_12433_0 & _T_16262;
  assign _GEN_465 = 5'h1 == _T_12733_0 ? _T_12514_0_1 : _T_12514_0_0;
  assign _GEN_466 = 5'h2 == _T_12733_0 ? _T_12514_0_2 : _GEN_465;
  assign _GEN_467 = 5'h3 == _T_12733_0 ? _T_12514_0_3 : _GEN_466;
  assign _GEN_468 = 5'h4 == _T_12733_0 ? _T_12514_0_4 : _GEN_467;
  assign _GEN_469 = 5'h5 == _T_12733_0 ? _T_12514_0_5 : _GEN_468;
  assign _GEN_470 = 5'h6 == _T_12733_0 ? _T_12514_0_6 : _GEN_469;
  assign _GEN_471 = 5'h7 == _T_12733_0 ? _T_12514_0_7 : _GEN_470;
  assign _GEN_472 = 5'h8 == _T_12733_0 ? _T_12514_0_8 : _GEN_471;
  assign _GEN_473 = 5'h9 == _T_12733_0 ? _T_12514_0_9 : _GEN_472;
  assign _GEN_474 = 5'ha == _T_12733_0 ? _T_12514_0_10 : _GEN_473;
  assign _GEN_475 = 5'hb == _T_12733_0 ? _T_12514_0_11 : _GEN_474;
  assign _GEN_476 = 5'hc == _T_12733_0 ? _T_12514_0_12 : _GEN_475;
  assign _GEN_477 = 5'hd == _T_12733_0 ? _T_12514_0_13 : _GEN_476;
  assign _GEN_478 = 5'he == _T_12733_0 ? _T_12514_0_14 : _GEN_477;
  assign _GEN_479 = 5'hf == _T_12733_0 ? _T_12514_0_15 : _GEN_478;
  assign _GEN_480 = 5'h10 == _T_12733_0 ? _T_12514_0_16 : _GEN_479;
  assign _GEN_481 = 5'h11 == _T_12733_0 ? _T_12514_0_17 : _GEN_480;
  assign _GEN_482 = 5'h12 == _T_12733_0 ? _T_12514_0_18 : _GEN_481;
  assign _GEN_483 = 5'h13 == _T_12733_0 ? _T_12514_0_19 : _GEN_482;
  assign _GEN_484 = 5'h14 == _T_12733_0 ? _T_12514_0_20 : _GEN_483;
  assign _GEN_485 = 5'h15 == _T_12733_0 ? _T_12514_0_21 : _GEN_484;
  assign _GEN_486 = 5'h16 == _T_12733_0 ? _T_12514_0_22 : _GEN_485;
  assign _GEN_487 = 5'h17 == _T_12733_0 ? _T_12514_0_23 : _GEN_486;
  assign _GEN_488 = 5'h18 == _T_12733_0 ? _T_12514_0_24 : _GEN_487;
  assign _GEN_489 = 5'h19 == _T_12733_0 ? _T_12514_0_25 : _GEN_488;
  assign _GEN_490 = 5'h1a == _T_12733_0 ? _T_12514_0_26 : _GEN_489;
  assign _GEN_491 = 5'h1b == _T_12733_0 ? _T_12514_0_27 : _GEN_490;
  assign _GEN_492 = 5'h1c == _T_12733_0 ? _T_12514_0_28 : _GEN_491;
  assign _GEN_493 = 5'h1d == _T_12733_0 ? _T_12514_0_29 : _GEN_492;
  assign _GEN_494 = 5'h1e == _T_12733_0 ? _T_12514_0_30 : _GEN_493;
  assign _GEN_495 = 5'h1f == _T_12733_0 ? _T_12514_0_31 : _GEN_494;
  assign _T_16305 = _T_407 - 1'h1;
  assign _T_16306 = $unsigned(_T_16305);
  assign _T_16307 = _T_16306[0:0];
  assign _T_16308 = _T_16278 ? 1'h0 : _T_16307;
  assign _T_16310 = 1'h0 < _T_12767;
  assign _T_16311 = _T_16310 ? _T_407 : _T_16308;
  assign _T_16313 = _T_16311 == 1'h0;
  assign _T_16315 = _T_16313 ? _T_12754_0 : 1'h0;
  assign _T_16322 = _T_16318 + 1'h1;
  assign _T_16323 = _T_16322[0:0];
  assign _GEN_496 = _T_16318 ? _T_16323 : _T_16318;
  assign _T_16346 = _T_16337_0 == 1'h0;
  assign _T_16670 = _T_16318 == 1'h0;
  assign _T_16672 = _T_16668 == 1'h0;
  assign _T_16673 = _T_16670 & _T_16672;
  assign _GEN_497 = _T_16673 ? 1'h1 : _T_16668;
  assign _T_16677 = _T_16670 & _T_506_0;
  assign _T_16679 = _T_518_0 == 5'h1f;
  assign _T_16680 = _T_16677 & _T_16679;
  assign _GEN_498 = _T_16680 ? 1'h1 : _T_16646_0;
  assign _GEN_499 = 5'h0 == _T_518_0 ? _GEN_4 : _T_16427_0_0;
  assign _GEN_500 = 5'h1 == _T_518_0 ? _GEN_4 : _T_16427_0_1;
  assign _GEN_501 = 5'h2 == _T_518_0 ? _GEN_4 : _T_16427_0_2;
  assign _GEN_502 = 5'h3 == _T_518_0 ? _GEN_4 : _T_16427_0_3;
  assign _GEN_503 = 5'h4 == _T_518_0 ? _GEN_4 : _T_16427_0_4;
  assign _GEN_504 = 5'h5 == _T_518_0 ? _GEN_4 : _T_16427_0_5;
  assign _GEN_505 = 5'h6 == _T_518_0 ? _GEN_4 : _T_16427_0_6;
  assign _GEN_506 = 5'h7 == _T_518_0 ? _GEN_4 : _T_16427_0_7;
  assign _GEN_507 = 5'h8 == _T_518_0 ? _GEN_4 : _T_16427_0_8;
  assign _GEN_508 = 5'h9 == _T_518_0 ? _GEN_4 : _T_16427_0_9;
  assign _GEN_509 = 5'ha == _T_518_0 ? _GEN_4 : _T_16427_0_10;
  assign _GEN_510 = 5'hb == _T_518_0 ? _GEN_4 : _T_16427_0_11;
  assign _GEN_511 = 5'hc == _T_518_0 ? _GEN_4 : _T_16427_0_12;
  assign _GEN_512 = 5'hd == _T_518_0 ? _GEN_4 : _T_16427_0_13;
  assign _GEN_513 = 5'he == _T_518_0 ? _GEN_4 : _T_16427_0_14;
  assign _GEN_514 = 5'hf == _T_518_0 ? _GEN_4 : _T_16427_0_15;
  assign _GEN_515 = 5'h10 == _T_518_0 ? _GEN_4 : _T_16427_0_16;
  assign _GEN_516 = 5'h11 == _T_518_0 ? _GEN_4 : _T_16427_0_17;
  assign _GEN_517 = 5'h12 == _T_518_0 ? _GEN_4 : _T_16427_0_18;
  assign _GEN_518 = 5'h13 == _T_518_0 ? _GEN_4 : _T_16427_0_19;
  assign _GEN_519 = 5'h14 == _T_518_0 ? _GEN_4 : _T_16427_0_20;
  assign _GEN_520 = 5'h15 == _T_518_0 ? _GEN_4 : _T_16427_0_21;
  assign _GEN_521 = 5'h16 == _T_518_0 ? _GEN_4 : _T_16427_0_22;
  assign _GEN_522 = 5'h17 == _T_518_0 ? _GEN_4 : _T_16427_0_23;
  assign _GEN_523 = 5'h18 == _T_518_0 ? _GEN_4 : _T_16427_0_24;
  assign _GEN_524 = 5'h19 == _T_518_0 ? _GEN_4 : _T_16427_0_25;
  assign _GEN_525 = 5'h1a == _T_518_0 ? _GEN_4 : _T_16427_0_26;
  assign _GEN_526 = 5'h1b == _T_518_0 ? _GEN_4 : _T_16427_0_27;
  assign _GEN_527 = 5'h1c == _T_518_0 ? _GEN_4 : _T_16427_0_28;
  assign _GEN_528 = 5'h1d == _T_518_0 ? _GEN_4 : _T_16427_0_29;
  assign _GEN_529 = 5'h1e == _T_518_0 ? _GEN_4 : _T_16427_0_30;
  assign _GEN_530 = 5'h1f == _T_518_0 ? _GEN_4 : _T_16427_0_31;
  assign _GEN_531 = _T_506_0 ? _GEN_499 : _T_16427_0_0;
  assign _GEN_532 = _T_506_0 ? _GEN_500 : _T_16427_0_1;
  assign _GEN_533 = _T_506_0 ? _GEN_501 : _T_16427_0_2;
  assign _GEN_534 = _T_506_0 ? _GEN_502 : _T_16427_0_3;
  assign _GEN_535 = _T_506_0 ? _GEN_503 : _T_16427_0_4;
  assign _GEN_536 = _T_506_0 ? _GEN_504 : _T_16427_0_5;
  assign _GEN_537 = _T_506_0 ? _GEN_505 : _T_16427_0_6;
  assign _GEN_538 = _T_506_0 ? _GEN_506 : _T_16427_0_7;
  assign _GEN_539 = _T_506_0 ? _GEN_507 : _T_16427_0_8;
  assign _GEN_540 = _T_506_0 ? _GEN_508 : _T_16427_0_9;
  assign _GEN_541 = _T_506_0 ? _GEN_509 : _T_16427_0_10;
  assign _GEN_542 = _T_506_0 ? _GEN_510 : _T_16427_0_11;
  assign _GEN_543 = _T_506_0 ? _GEN_511 : _T_16427_0_12;
  assign _GEN_544 = _T_506_0 ? _GEN_512 : _T_16427_0_13;
  assign _GEN_545 = _T_506_0 ? _GEN_513 : _T_16427_0_14;
  assign _GEN_546 = _T_506_0 ? _GEN_514 : _T_16427_0_15;
  assign _GEN_547 = _T_506_0 ? _GEN_515 : _T_16427_0_16;
  assign _GEN_548 = _T_506_0 ? _GEN_516 : _T_16427_0_17;
  assign _GEN_549 = _T_506_0 ? _GEN_517 : _T_16427_0_18;
  assign _GEN_550 = _T_506_0 ? _GEN_518 : _T_16427_0_19;
  assign _GEN_551 = _T_506_0 ? _GEN_519 : _T_16427_0_20;
  assign _GEN_552 = _T_506_0 ? _GEN_520 : _T_16427_0_21;
  assign _GEN_553 = _T_506_0 ? _GEN_521 : _T_16427_0_22;
  assign _GEN_554 = _T_506_0 ? _GEN_522 : _T_16427_0_23;
  assign _GEN_555 = _T_506_0 ? _GEN_523 : _T_16427_0_24;
  assign _GEN_556 = _T_506_0 ? _GEN_524 : _T_16427_0_25;
  assign _GEN_557 = _T_506_0 ? _GEN_525 : _T_16427_0_26;
  assign _GEN_558 = _T_506_0 ? _GEN_526 : _T_16427_0_27;
  assign _GEN_559 = _T_506_0 ? _GEN_527 : _T_16427_0_28;
  assign _GEN_560 = _T_506_0 ? _GEN_528 : _T_16427_0_29;
  assign _GEN_561 = _T_506_0 ? _GEN_529 : _T_16427_0_30;
  assign _GEN_562 = _T_506_0 ? _GEN_530 : _T_16427_0_31;
  assign _T_16686 = _T_16670 & _T_500_0;
  assign _T_16689 = _T_16686 & _T_16346;
  assign _T_16695 = _T_16689 & _T_16672;
  assign _GEN_563 = _T_16695 ? 1'h1 : _T_16337_0;
  assign _GEN_564 = _T_16695 ? _T_494_0 : _T_16350_0;
  assign _T_16704 = _T_16659 == 1'h0;
  assign _T_16705 = _T_16337_0 & _T_16704;
  assign _T_16810 = {_T_16427_0_1,_T_16427_0_0};
  assign _T_16811 = {_T_16427_0_3,_T_16427_0_2};
  assign _T_16812 = {_T_16811,_T_16810};
  assign _T_16813 = {_T_16427_0_5,_T_16427_0_4};
  assign _T_16814 = {_T_16427_0_7,_T_16427_0_6};
  assign _T_16815 = {_T_16814,_T_16813};
  assign _T_16816 = {_T_16815,_T_16812};
  assign _T_16817 = {_T_16427_0_9,_T_16427_0_8};
  assign _T_16818 = {_T_16427_0_11,_T_16427_0_10};
  assign _T_16819 = {_T_16818,_T_16817};
  assign _T_16820 = {_T_16427_0_13,_T_16427_0_12};
  assign _T_16821 = {_T_16427_0_15,_T_16427_0_14};
  assign _T_16822 = {_T_16821,_T_16820};
  assign _T_16823 = {_T_16822,_T_16819};
  assign _T_16824 = {_T_16823,_T_16816};
  assign _T_16825 = {_T_16427_0_17,_T_16427_0_16};
  assign _T_16826 = {_T_16427_0_19,_T_16427_0_18};
  assign _T_16827 = {_T_16826,_T_16825};
  assign _T_16828 = {_T_16427_0_21,_T_16427_0_20};
  assign _T_16829 = {_T_16427_0_23,_T_16427_0_22};
  assign _T_16830 = {_T_16829,_T_16828};
  assign _T_16831 = {_T_16830,_T_16827};
  assign _T_16832 = {_T_16427_0_25,_T_16427_0_24};
  assign _T_16833 = {_T_16427_0_27,_T_16427_0_26};
  assign _T_16834 = {_T_16833,_T_16832};
  assign _T_16835 = {_T_16427_0_29,_T_16427_0_28};
  assign _T_16836 = {_T_16427_0_31,_T_16427_0_30};
  assign _T_16837 = {_T_16836,_T_16835};
  assign _T_16838 = {_T_16837,_T_16834};
  assign _T_16839 = {_T_16838,_T_16831};
  assign _T_16840 = {_T_16839,_T_16824};
  assign _T_16841 = _T_16840[511:0];
  assign _T_16844 = _T_16840[1023:512];
  assign _T_16845 = _T_16665 ? _T_16844 : _T_16841;
  assign _T_16852 = io_axi_outputMemAddrValids_0 & io_axi_outputMemAddrReadys_0;
  assign _T_16859 = _T_16668 & _T_16346;
  assign _T_16860 = _T_16852 | _T_16859;
  assign _T_16862 = _T_16656 == 1'h0;
  assign _T_16865 = _T_16656 + 1'h1;
  assign _T_16866 = _T_16865[0:0];
  assign _GEN_565 = _T_16862 ? 1'h1 : _T_16659;
  assign _GEN_566 = _T_16862 ? _T_16656 : _T_16866;
  assign _GEN_567 = _T_16860 ? _GEN_565 : _T_16659;
  assign _GEN_568 = _T_16860 ? _GEN_566 : _T_16656;
  assign _T_16867 = io_axi_outputMemBlockValids_0 & io_axi_outputMemBlockReadys_0;
  assign _T_16872 = _T_16665 + 1'h1;
  assign _T_16873 = _T_16872[0:0];
  assign _T_16874 = _T_16665 ? 1'h0 : _T_16873;
  assign _GEN_569 = _T_16867 ? _T_16874 : _T_16665;
  assign _T_16878 = _T_16867 & _T_16665;
  assign _T_16885 = _T_16662 < _T_16656;
  assign _T_16886 = _T_16885 | _T_16659;
  assign _T_16887 = _T_16346 & _T_16886;
  assign _T_16888 = _T_16878 | _T_16887;
  assign _T_16890 = _T_16662 == 1'h0;
  assign _T_16892 = _T_410 == 1'h0;
  assign _T_16895 = _T_410 + 1'h1;
  assign _T_16896 = _T_16895[0:0];
  assign _T_16897 = _T_16892 ? 1'h0 : _T_16896;
  assign _T_16906 = _T_16662 + 1'h1;
  assign _T_16907 = _T_16906[0:0];
  assign _GEN_570 = _T_16890 ? _T_16897 : _T_410;
  assign _GEN_571 = _T_16890 ? 1'h0 : _GEN_496;
  assign _GEN_572 = _T_16890 ? 1'h0 : _T_16907;
  assign _GEN_573 = _T_16890 ? 1'h0 : _GEN_568;
  assign _GEN_574 = _T_16890 ? 1'h0 : _GEN_567;
  assign _GEN_575 = _T_16890 ? 1'h0 : _GEN_497;
  assign _GEN_576 = _T_16890 ? 1'h0 : _GEN_563;
  assign _GEN_577 = _T_16890 ? 1'h0 : _GEN_498;
  assign _GEN_578 = _T_16888 ? _GEN_570 : _T_410;
  assign _GEN_579 = _T_16888 ? _GEN_571 : _GEN_496;
  assign _GEN_580 = _T_16888 ? _GEN_572 : _T_16662;
  assign _GEN_581 = _T_16888 ? _GEN_573 : _GEN_568;
  assign _GEN_582 = _T_16888 ? _GEN_574 : _GEN_567;
  assign _GEN_583 = _T_16888 ? _GEN_575 : _GEN_497;
  assign _GEN_584 = _T_16888 ? _GEN_576 : _GEN_563;
  assign _GEN_585 = _T_16888 ? _GEN_577 : _GEN_498;
  assign _T_16923 = _T_16892 ? _T_16695 : 1'h0;
  assign _T_16930 = _T_16926 + 1'h1;
  assign _T_16931 = _T_16930[0:0];
  assign _GEN_586 = _T_16926 ? _T_16931 : _T_16926;
  assign _T_16954 = _T_16945_0 == 1'h0;
  assign _T_17278 = _T_16926 == 1'h0;
  assign _T_17280 = _T_17276 == 1'h0;
  assign _T_17281 = _T_17278 & _T_17280;
  assign _GEN_587 = _T_17281 ? 1'h1 : _T_17276;
  assign _T_17285 = _T_17278 & _T_542_0;
  assign _T_17287 = _T_554_0 == 5'h1f;
  assign _T_17288 = _T_17285 & _T_17287;
  assign _GEN_588 = _T_17288 ? 1'h1 : _T_17254_0;
  assign _GEN_589 = 5'h0 == _T_554_0 ? _GEN_5 : _T_17035_0_0;
  assign _GEN_590 = 5'h1 == _T_554_0 ? _GEN_5 : _T_17035_0_1;
  assign _GEN_591 = 5'h2 == _T_554_0 ? _GEN_5 : _T_17035_0_2;
  assign _GEN_592 = 5'h3 == _T_554_0 ? _GEN_5 : _T_17035_0_3;
  assign _GEN_593 = 5'h4 == _T_554_0 ? _GEN_5 : _T_17035_0_4;
  assign _GEN_594 = 5'h5 == _T_554_0 ? _GEN_5 : _T_17035_0_5;
  assign _GEN_595 = 5'h6 == _T_554_0 ? _GEN_5 : _T_17035_0_6;
  assign _GEN_596 = 5'h7 == _T_554_0 ? _GEN_5 : _T_17035_0_7;
  assign _GEN_597 = 5'h8 == _T_554_0 ? _GEN_5 : _T_17035_0_8;
  assign _GEN_598 = 5'h9 == _T_554_0 ? _GEN_5 : _T_17035_0_9;
  assign _GEN_599 = 5'ha == _T_554_0 ? _GEN_5 : _T_17035_0_10;
  assign _GEN_600 = 5'hb == _T_554_0 ? _GEN_5 : _T_17035_0_11;
  assign _GEN_601 = 5'hc == _T_554_0 ? _GEN_5 : _T_17035_0_12;
  assign _GEN_602 = 5'hd == _T_554_0 ? _GEN_5 : _T_17035_0_13;
  assign _GEN_603 = 5'he == _T_554_0 ? _GEN_5 : _T_17035_0_14;
  assign _GEN_604 = 5'hf == _T_554_0 ? _GEN_5 : _T_17035_0_15;
  assign _GEN_605 = 5'h10 == _T_554_0 ? _GEN_5 : _T_17035_0_16;
  assign _GEN_606 = 5'h11 == _T_554_0 ? _GEN_5 : _T_17035_0_17;
  assign _GEN_607 = 5'h12 == _T_554_0 ? _GEN_5 : _T_17035_0_18;
  assign _GEN_608 = 5'h13 == _T_554_0 ? _GEN_5 : _T_17035_0_19;
  assign _GEN_609 = 5'h14 == _T_554_0 ? _GEN_5 : _T_17035_0_20;
  assign _GEN_610 = 5'h15 == _T_554_0 ? _GEN_5 : _T_17035_0_21;
  assign _GEN_611 = 5'h16 == _T_554_0 ? _GEN_5 : _T_17035_0_22;
  assign _GEN_612 = 5'h17 == _T_554_0 ? _GEN_5 : _T_17035_0_23;
  assign _GEN_613 = 5'h18 == _T_554_0 ? _GEN_5 : _T_17035_0_24;
  assign _GEN_614 = 5'h19 == _T_554_0 ? _GEN_5 : _T_17035_0_25;
  assign _GEN_615 = 5'h1a == _T_554_0 ? _GEN_5 : _T_17035_0_26;
  assign _GEN_616 = 5'h1b == _T_554_0 ? _GEN_5 : _T_17035_0_27;
  assign _GEN_617 = 5'h1c == _T_554_0 ? _GEN_5 : _T_17035_0_28;
  assign _GEN_618 = 5'h1d == _T_554_0 ? _GEN_5 : _T_17035_0_29;
  assign _GEN_619 = 5'h1e == _T_554_0 ? _GEN_5 : _T_17035_0_30;
  assign _GEN_620 = 5'h1f == _T_554_0 ? _GEN_5 : _T_17035_0_31;
  assign _GEN_621 = _T_542_0 ? _GEN_589 : _T_17035_0_0;
  assign _GEN_622 = _T_542_0 ? _GEN_590 : _T_17035_0_1;
  assign _GEN_623 = _T_542_0 ? _GEN_591 : _T_17035_0_2;
  assign _GEN_624 = _T_542_0 ? _GEN_592 : _T_17035_0_3;
  assign _GEN_625 = _T_542_0 ? _GEN_593 : _T_17035_0_4;
  assign _GEN_626 = _T_542_0 ? _GEN_594 : _T_17035_0_5;
  assign _GEN_627 = _T_542_0 ? _GEN_595 : _T_17035_0_6;
  assign _GEN_628 = _T_542_0 ? _GEN_596 : _T_17035_0_7;
  assign _GEN_629 = _T_542_0 ? _GEN_597 : _T_17035_0_8;
  assign _GEN_630 = _T_542_0 ? _GEN_598 : _T_17035_0_9;
  assign _GEN_631 = _T_542_0 ? _GEN_599 : _T_17035_0_10;
  assign _GEN_632 = _T_542_0 ? _GEN_600 : _T_17035_0_11;
  assign _GEN_633 = _T_542_0 ? _GEN_601 : _T_17035_0_12;
  assign _GEN_634 = _T_542_0 ? _GEN_602 : _T_17035_0_13;
  assign _GEN_635 = _T_542_0 ? _GEN_603 : _T_17035_0_14;
  assign _GEN_636 = _T_542_0 ? _GEN_604 : _T_17035_0_15;
  assign _GEN_637 = _T_542_0 ? _GEN_605 : _T_17035_0_16;
  assign _GEN_638 = _T_542_0 ? _GEN_606 : _T_17035_0_17;
  assign _GEN_639 = _T_542_0 ? _GEN_607 : _T_17035_0_18;
  assign _GEN_640 = _T_542_0 ? _GEN_608 : _T_17035_0_19;
  assign _GEN_641 = _T_542_0 ? _GEN_609 : _T_17035_0_20;
  assign _GEN_642 = _T_542_0 ? _GEN_610 : _T_17035_0_21;
  assign _GEN_643 = _T_542_0 ? _GEN_611 : _T_17035_0_22;
  assign _GEN_644 = _T_542_0 ? _GEN_612 : _T_17035_0_23;
  assign _GEN_645 = _T_542_0 ? _GEN_613 : _T_17035_0_24;
  assign _GEN_646 = _T_542_0 ? _GEN_614 : _T_17035_0_25;
  assign _GEN_647 = _T_542_0 ? _GEN_615 : _T_17035_0_26;
  assign _GEN_648 = _T_542_0 ? _GEN_616 : _T_17035_0_27;
  assign _GEN_649 = _T_542_0 ? _GEN_617 : _T_17035_0_28;
  assign _GEN_650 = _T_542_0 ? _GEN_618 : _T_17035_0_29;
  assign _GEN_651 = _T_542_0 ? _GEN_619 : _T_17035_0_30;
  assign _GEN_652 = _T_542_0 ? _GEN_620 : _T_17035_0_31;
  assign _T_17294 = _T_17278 & _T_536_0;
  assign _T_17297 = _T_17294 & _T_16954;
  assign _T_17303 = _T_17297 & _T_17280;
  assign _GEN_653 = _T_17303 ? 1'h1 : _T_16945_0;
  assign _GEN_654 = _T_17303 ? _T_530_0 : _T_16958_0;
  assign _T_17312 = _T_17267 == 1'h0;
  assign _T_17313 = _T_16945_0 & _T_17312;
  assign _T_17418 = {_T_17035_0_1,_T_17035_0_0};
  assign _T_17419 = {_T_17035_0_3,_T_17035_0_2};
  assign _T_17420 = {_T_17419,_T_17418};
  assign _T_17421 = {_T_17035_0_5,_T_17035_0_4};
  assign _T_17422 = {_T_17035_0_7,_T_17035_0_6};
  assign _T_17423 = {_T_17422,_T_17421};
  assign _T_17424 = {_T_17423,_T_17420};
  assign _T_17425 = {_T_17035_0_9,_T_17035_0_8};
  assign _T_17426 = {_T_17035_0_11,_T_17035_0_10};
  assign _T_17427 = {_T_17426,_T_17425};
  assign _T_17428 = {_T_17035_0_13,_T_17035_0_12};
  assign _T_17429 = {_T_17035_0_15,_T_17035_0_14};
  assign _T_17430 = {_T_17429,_T_17428};
  assign _T_17431 = {_T_17430,_T_17427};
  assign _T_17432 = {_T_17431,_T_17424};
  assign _T_17433 = {_T_17035_0_17,_T_17035_0_16};
  assign _T_17434 = {_T_17035_0_19,_T_17035_0_18};
  assign _T_17435 = {_T_17434,_T_17433};
  assign _T_17436 = {_T_17035_0_21,_T_17035_0_20};
  assign _T_17437 = {_T_17035_0_23,_T_17035_0_22};
  assign _T_17438 = {_T_17437,_T_17436};
  assign _T_17439 = {_T_17438,_T_17435};
  assign _T_17440 = {_T_17035_0_25,_T_17035_0_24};
  assign _T_17441 = {_T_17035_0_27,_T_17035_0_26};
  assign _T_17442 = {_T_17441,_T_17440};
  assign _T_17443 = {_T_17035_0_29,_T_17035_0_28};
  assign _T_17444 = {_T_17035_0_31,_T_17035_0_30};
  assign _T_17445 = {_T_17444,_T_17443};
  assign _T_17446 = {_T_17445,_T_17442};
  assign _T_17447 = {_T_17446,_T_17439};
  assign _T_17448 = {_T_17447,_T_17432};
  assign _T_17449 = _T_17448[511:0];
  assign _T_17452 = _T_17448[1023:512];
  assign _T_17453 = _T_17273 ? _T_17452 : _T_17449;
  assign _T_17460 = io_axi_outputMemAddrValids_1 & io_axi_outputMemAddrReadys_1;
  assign _T_17467 = _T_17276 & _T_16954;
  assign _T_17468 = _T_17460 | _T_17467;
  assign _T_17470 = _T_17264 == 1'h0;
  assign _T_17473 = _T_17264 + 1'h1;
  assign _T_17474 = _T_17473[0:0];
  assign _GEN_655 = _T_17470 ? 1'h1 : _T_17267;
  assign _GEN_656 = _T_17470 ? _T_17264 : _T_17474;
  assign _GEN_657 = _T_17468 ? _GEN_655 : _T_17267;
  assign _GEN_658 = _T_17468 ? _GEN_656 : _T_17264;
  assign _T_17475 = io_axi_outputMemBlockValids_1 & io_axi_outputMemBlockReadys_1;
  assign _T_17480 = _T_17273 + 1'h1;
  assign _T_17481 = _T_17480[0:0];
  assign _T_17482 = _T_17273 ? 1'h0 : _T_17481;
  assign _GEN_659 = _T_17475 ? _T_17482 : _T_17273;
  assign _T_17486 = _T_17475 & _T_17273;
  assign _T_17493 = _T_17270 < _T_17264;
  assign _T_17494 = _T_17493 | _T_17267;
  assign _T_17495 = _T_16954 & _T_17494;
  assign _T_17496 = _T_17486 | _T_17495;
  assign _T_17498 = _T_17270 == 1'h0;
  assign _T_17500 = _T_413 == 1'h0;
  assign _T_17503 = _T_413 + 1'h1;
  assign _T_17504 = _T_17503[0:0];
  assign _T_17505 = _T_17500 ? 1'h0 : _T_17504;
  assign _T_17514 = _T_17270 + 1'h1;
  assign _T_17515 = _T_17514[0:0];
  assign _GEN_660 = _T_17498 ? _T_17505 : _T_413;
  assign _GEN_661 = _T_17498 ? 1'h0 : _GEN_586;
  assign _GEN_662 = _T_17498 ? 1'h0 : _T_17515;
  assign _GEN_663 = _T_17498 ? 1'h0 : _GEN_658;
  assign _GEN_664 = _T_17498 ? 1'h0 : _GEN_657;
  assign _GEN_665 = _T_17498 ? 1'h0 : _GEN_587;
  assign _GEN_666 = _T_17498 ? 1'h0 : _GEN_653;
  assign _GEN_667 = _T_17498 ? 1'h0 : _GEN_588;
  assign _GEN_668 = _T_17496 ? _GEN_660 : _T_413;
  assign _GEN_669 = _T_17496 ? _GEN_661 : _GEN_586;
  assign _GEN_670 = _T_17496 ? _GEN_662 : _T_17270;
  assign _GEN_671 = _T_17496 ? _GEN_663 : _GEN_658;
  assign _GEN_672 = _T_17496 ? _GEN_664 : _GEN_657;
  assign _GEN_673 = _T_17496 ? _GEN_665 : _GEN_587;
  assign _GEN_674 = _T_17496 ? _GEN_666 : _GEN_653;
  assign _GEN_675 = _T_17496 ? _GEN_667 : _GEN_588;
  assign _T_17531 = _T_17500 ? _T_17303 : 1'h0;
  assign _T_17538 = _T_17534 + 1'h1;
  assign _T_17539 = _T_17538[0:0];
  assign _GEN_676 = _T_17534 ? _T_17539 : _T_17534;
  assign _T_17562 = _T_17553_0 == 1'h0;
  assign _T_17886 = _T_17534 == 1'h0;
  assign _T_17888 = _T_17884 == 1'h0;
  assign _T_17889 = _T_17886 & _T_17888;
  assign _GEN_677 = _T_17889 ? 1'h1 : _T_17884;
  assign _T_17893 = _T_17886 & _T_578_0;
  assign _T_17895 = _T_590_0 == 5'h1f;
  assign _T_17896 = _T_17893 & _T_17895;
  assign _GEN_678 = _T_17896 ? 1'h1 : _T_17862_0;
  assign _GEN_679 = 5'h0 == _T_590_0 ? _GEN_6 : _T_17643_0_0;
  assign _GEN_680 = 5'h1 == _T_590_0 ? _GEN_6 : _T_17643_0_1;
  assign _GEN_681 = 5'h2 == _T_590_0 ? _GEN_6 : _T_17643_0_2;
  assign _GEN_682 = 5'h3 == _T_590_0 ? _GEN_6 : _T_17643_0_3;
  assign _GEN_683 = 5'h4 == _T_590_0 ? _GEN_6 : _T_17643_0_4;
  assign _GEN_684 = 5'h5 == _T_590_0 ? _GEN_6 : _T_17643_0_5;
  assign _GEN_685 = 5'h6 == _T_590_0 ? _GEN_6 : _T_17643_0_6;
  assign _GEN_686 = 5'h7 == _T_590_0 ? _GEN_6 : _T_17643_0_7;
  assign _GEN_687 = 5'h8 == _T_590_0 ? _GEN_6 : _T_17643_0_8;
  assign _GEN_688 = 5'h9 == _T_590_0 ? _GEN_6 : _T_17643_0_9;
  assign _GEN_689 = 5'ha == _T_590_0 ? _GEN_6 : _T_17643_0_10;
  assign _GEN_690 = 5'hb == _T_590_0 ? _GEN_6 : _T_17643_0_11;
  assign _GEN_691 = 5'hc == _T_590_0 ? _GEN_6 : _T_17643_0_12;
  assign _GEN_692 = 5'hd == _T_590_0 ? _GEN_6 : _T_17643_0_13;
  assign _GEN_693 = 5'he == _T_590_0 ? _GEN_6 : _T_17643_0_14;
  assign _GEN_694 = 5'hf == _T_590_0 ? _GEN_6 : _T_17643_0_15;
  assign _GEN_695 = 5'h10 == _T_590_0 ? _GEN_6 : _T_17643_0_16;
  assign _GEN_696 = 5'h11 == _T_590_0 ? _GEN_6 : _T_17643_0_17;
  assign _GEN_697 = 5'h12 == _T_590_0 ? _GEN_6 : _T_17643_0_18;
  assign _GEN_698 = 5'h13 == _T_590_0 ? _GEN_6 : _T_17643_0_19;
  assign _GEN_699 = 5'h14 == _T_590_0 ? _GEN_6 : _T_17643_0_20;
  assign _GEN_700 = 5'h15 == _T_590_0 ? _GEN_6 : _T_17643_0_21;
  assign _GEN_701 = 5'h16 == _T_590_0 ? _GEN_6 : _T_17643_0_22;
  assign _GEN_702 = 5'h17 == _T_590_0 ? _GEN_6 : _T_17643_0_23;
  assign _GEN_703 = 5'h18 == _T_590_0 ? _GEN_6 : _T_17643_0_24;
  assign _GEN_704 = 5'h19 == _T_590_0 ? _GEN_6 : _T_17643_0_25;
  assign _GEN_705 = 5'h1a == _T_590_0 ? _GEN_6 : _T_17643_0_26;
  assign _GEN_706 = 5'h1b == _T_590_0 ? _GEN_6 : _T_17643_0_27;
  assign _GEN_707 = 5'h1c == _T_590_0 ? _GEN_6 : _T_17643_0_28;
  assign _GEN_708 = 5'h1d == _T_590_0 ? _GEN_6 : _T_17643_0_29;
  assign _GEN_709 = 5'h1e == _T_590_0 ? _GEN_6 : _T_17643_0_30;
  assign _GEN_710 = 5'h1f == _T_590_0 ? _GEN_6 : _T_17643_0_31;
  assign _GEN_711 = _T_578_0 ? _GEN_679 : _T_17643_0_0;
  assign _GEN_712 = _T_578_0 ? _GEN_680 : _T_17643_0_1;
  assign _GEN_713 = _T_578_0 ? _GEN_681 : _T_17643_0_2;
  assign _GEN_714 = _T_578_0 ? _GEN_682 : _T_17643_0_3;
  assign _GEN_715 = _T_578_0 ? _GEN_683 : _T_17643_0_4;
  assign _GEN_716 = _T_578_0 ? _GEN_684 : _T_17643_0_5;
  assign _GEN_717 = _T_578_0 ? _GEN_685 : _T_17643_0_6;
  assign _GEN_718 = _T_578_0 ? _GEN_686 : _T_17643_0_7;
  assign _GEN_719 = _T_578_0 ? _GEN_687 : _T_17643_0_8;
  assign _GEN_720 = _T_578_0 ? _GEN_688 : _T_17643_0_9;
  assign _GEN_721 = _T_578_0 ? _GEN_689 : _T_17643_0_10;
  assign _GEN_722 = _T_578_0 ? _GEN_690 : _T_17643_0_11;
  assign _GEN_723 = _T_578_0 ? _GEN_691 : _T_17643_0_12;
  assign _GEN_724 = _T_578_0 ? _GEN_692 : _T_17643_0_13;
  assign _GEN_725 = _T_578_0 ? _GEN_693 : _T_17643_0_14;
  assign _GEN_726 = _T_578_0 ? _GEN_694 : _T_17643_0_15;
  assign _GEN_727 = _T_578_0 ? _GEN_695 : _T_17643_0_16;
  assign _GEN_728 = _T_578_0 ? _GEN_696 : _T_17643_0_17;
  assign _GEN_729 = _T_578_0 ? _GEN_697 : _T_17643_0_18;
  assign _GEN_730 = _T_578_0 ? _GEN_698 : _T_17643_0_19;
  assign _GEN_731 = _T_578_0 ? _GEN_699 : _T_17643_0_20;
  assign _GEN_732 = _T_578_0 ? _GEN_700 : _T_17643_0_21;
  assign _GEN_733 = _T_578_0 ? _GEN_701 : _T_17643_0_22;
  assign _GEN_734 = _T_578_0 ? _GEN_702 : _T_17643_0_23;
  assign _GEN_735 = _T_578_0 ? _GEN_703 : _T_17643_0_24;
  assign _GEN_736 = _T_578_0 ? _GEN_704 : _T_17643_0_25;
  assign _GEN_737 = _T_578_0 ? _GEN_705 : _T_17643_0_26;
  assign _GEN_738 = _T_578_0 ? _GEN_706 : _T_17643_0_27;
  assign _GEN_739 = _T_578_0 ? _GEN_707 : _T_17643_0_28;
  assign _GEN_740 = _T_578_0 ? _GEN_708 : _T_17643_0_29;
  assign _GEN_741 = _T_578_0 ? _GEN_709 : _T_17643_0_30;
  assign _GEN_742 = _T_578_0 ? _GEN_710 : _T_17643_0_31;
  assign _T_17902 = _T_17886 & _T_572_0;
  assign _T_17905 = _T_17902 & _T_17562;
  assign _T_17911 = _T_17905 & _T_17888;
  assign _GEN_743 = _T_17911 ? 1'h1 : _T_17553_0;
  assign _GEN_744 = _T_17911 ? _T_566_0 : _T_17566_0;
  assign _T_17920 = _T_17875 == 1'h0;
  assign _T_17921 = _T_17553_0 & _T_17920;
  assign _T_18026 = {_T_17643_0_1,_T_17643_0_0};
  assign _T_18027 = {_T_17643_0_3,_T_17643_0_2};
  assign _T_18028 = {_T_18027,_T_18026};
  assign _T_18029 = {_T_17643_0_5,_T_17643_0_4};
  assign _T_18030 = {_T_17643_0_7,_T_17643_0_6};
  assign _T_18031 = {_T_18030,_T_18029};
  assign _T_18032 = {_T_18031,_T_18028};
  assign _T_18033 = {_T_17643_0_9,_T_17643_0_8};
  assign _T_18034 = {_T_17643_0_11,_T_17643_0_10};
  assign _T_18035 = {_T_18034,_T_18033};
  assign _T_18036 = {_T_17643_0_13,_T_17643_0_12};
  assign _T_18037 = {_T_17643_0_15,_T_17643_0_14};
  assign _T_18038 = {_T_18037,_T_18036};
  assign _T_18039 = {_T_18038,_T_18035};
  assign _T_18040 = {_T_18039,_T_18032};
  assign _T_18041 = {_T_17643_0_17,_T_17643_0_16};
  assign _T_18042 = {_T_17643_0_19,_T_17643_0_18};
  assign _T_18043 = {_T_18042,_T_18041};
  assign _T_18044 = {_T_17643_0_21,_T_17643_0_20};
  assign _T_18045 = {_T_17643_0_23,_T_17643_0_22};
  assign _T_18046 = {_T_18045,_T_18044};
  assign _T_18047 = {_T_18046,_T_18043};
  assign _T_18048 = {_T_17643_0_25,_T_17643_0_24};
  assign _T_18049 = {_T_17643_0_27,_T_17643_0_26};
  assign _T_18050 = {_T_18049,_T_18048};
  assign _T_18051 = {_T_17643_0_29,_T_17643_0_28};
  assign _T_18052 = {_T_17643_0_31,_T_17643_0_30};
  assign _T_18053 = {_T_18052,_T_18051};
  assign _T_18054 = {_T_18053,_T_18050};
  assign _T_18055 = {_T_18054,_T_18047};
  assign _T_18056 = {_T_18055,_T_18040};
  assign _T_18057 = _T_18056[511:0];
  assign _T_18060 = _T_18056[1023:512];
  assign _T_18061 = _T_17881 ? _T_18060 : _T_18057;
  assign _T_18068 = io_axi_outputMemAddrValids_2 & io_axi_outputMemAddrReadys_2;
  assign _T_18075 = _T_17884 & _T_17562;
  assign _T_18076 = _T_18068 | _T_18075;
  assign _T_18078 = _T_17872 == 1'h0;
  assign _T_18081 = _T_17872 + 1'h1;
  assign _T_18082 = _T_18081[0:0];
  assign _GEN_745 = _T_18078 ? 1'h1 : _T_17875;
  assign _GEN_746 = _T_18078 ? _T_17872 : _T_18082;
  assign _GEN_747 = _T_18076 ? _GEN_745 : _T_17875;
  assign _GEN_748 = _T_18076 ? _GEN_746 : _T_17872;
  assign _T_18083 = io_axi_outputMemBlockValids_2 & io_axi_outputMemBlockReadys_2;
  assign _T_18088 = _T_17881 + 1'h1;
  assign _T_18089 = _T_18088[0:0];
  assign _T_18090 = _T_17881 ? 1'h0 : _T_18089;
  assign _GEN_749 = _T_18083 ? _T_18090 : _T_17881;
  assign _T_18094 = _T_18083 & _T_17881;
  assign _T_18101 = _T_17878 < _T_17872;
  assign _T_18102 = _T_18101 | _T_17875;
  assign _T_18103 = _T_17562 & _T_18102;
  assign _T_18104 = _T_18094 | _T_18103;
  assign _T_18106 = _T_17878 == 1'h0;
  assign _T_18108 = _T_416 == 1'h0;
  assign _T_18111 = _T_416 + 1'h1;
  assign _T_18112 = _T_18111[0:0];
  assign _T_18113 = _T_18108 ? 1'h0 : _T_18112;
  assign _T_18122 = _T_17878 + 1'h1;
  assign _T_18123 = _T_18122[0:0];
  assign _GEN_750 = _T_18106 ? _T_18113 : _T_416;
  assign _GEN_751 = _T_18106 ? 1'h0 : _GEN_676;
  assign _GEN_752 = _T_18106 ? 1'h0 : _T_18123;
  assign _GEN_753 = _T_18106 ? 1'h0 : _GEN_748;
  assign _GEN_754 = _T_18106 ? 1'h0 : _GEN_747;
  assign _GEN_755 = _T_18106 ? 1'h0 : _GEN_677;
  assign _GEN_756 = _T_18106 ? 1'h0 : _GEN_743;
  assign _GEN_757 = _T_18106 ? 1'h0 : _GEN_678;
  assign _GEN_758 = _T_18104 ? _GEN_750 : _T_416;
  assign _GEN_759 = _T_18104 ? _GEN_751 : _GEN_676;
  assign _GEN_760 = _T_18104 ? _GEN_752 : _T_17878;
  assign _GEN_761 = _T_18104 ? _GEN_753 : _GEN_748;
  assign _GEN_762 = _T_18104 ? _GEN_754 : _GEN_747;
  assign _GEN_763 = _T_18104 ? _GEN_755 : _GEN_677;
  assign _GEN_764 = _T_18104 ? _GEN_756 : _GEN_743;
  assign _GEN_765 = _T_18104 ? _GEN_757 : _GEN_678;
  assign _T_18139 = _T_18108 ? _T_17911 : 1'h0;
  assign _T_18146 = _T_18142 + 1'h1;
  assign _T_18147 = _T_18146[0:0];
  assign _GEN_766 = _T_18142 ? _T_18147 : _T_18142;
  assign _T_18170 = _T_18161_0 == 1'h0;
  assign _T_18494 = _T_18142 == 1'h0;
  assign _T_18496 = _T_18492 == 1'h0;
  assign _T_18497 = _T_18494 & _T_18496;
  assign _GEN_767 = _T_18497 ? 1'h1 : _T_18492;
  assign _T_18501 = _T_18494 & _T_614_0;
  assign _T_18503 = _T_626_0 == 5'h1f;
  assign _T_18504 = _T_18501 & _T_18503;
  assign _GEN_768 = _T_18504 ? 1'h1 : _T_18470_0;
  assign _GEN_769 = 5'h0 == _T_626_0 ? _GEN_7 : _T_18251_0_0;
  assign _GEN_770 = 5'h1 == _T_626_0 ? _GEN_7 : _T_18251_0_1;
  assign _GEN_771 = 5'h2 == _T_626_0 ? _GEN_7 : _T_18251_0_2;
  assign _GEN_772 = 5'h3 == _T_626_0 ? _GEN_7 : _T_18251_0_3;
  assign _GEN_773 = 5'h4 == _T_626_0 ? _GEN_7 : _T_18251_0_4;
  assign _GEN_774 = 5'h5 == _T_626_0 ? _GEN_7 : _T_18251_0_5;
  assign _GEN_775 = 5'h6 == _T_626_0 ? _GEN_7 : _T_18251_0_6;
  assign _GEN_776 = 5'h7 == _T_626_0 ? _GEN_7 : _T_18251_0_7;
  assign _GEN_777 = 5'h8 == _T_626_0 ? _GEN_7 : _T_18251_0_8;
  assign _GEN_778 = 5'h9 == _T_626_0 ? _GEN_7 : _T_18251_0_9;
  assign _GEN_779 = 5'ha == _T_626_0 ? _GEN_7 : _T_18251_0_10;
  assign _GEN_780 = 5'hb == _T_626_0 ? _GEN_7 : _T_18251_0_11;
  assign _GEN_781 = 5'hc == _T_626_0 ? _GEN_7 : _T_18251_0_12;
  assign _GEN_782 = 5'hd == _T_626_0 ? _GEN_7 : _T_18251_0_13;
  assign _GEN_783 = 5'he == _T_626_0 ? _GEN_7 : _T_18251_0_14;
  assign _GEN_784 = 5'hf == _T_626_0 ? _GEN_7 : _T_18251_0_15;
  assign _GEN_785 = 5'h10 == _T_626_0 ? _GEN_7 : _T_18251_0_16;
  assign _GEN_786 = 5'h11 == _T_626_0 ? _GEN_7 : _T_18251_0_17;
  assign _GEN_787 = 5'h12 == _T_626_0 ? _GEN_7 : _T_18251_0_18;
  assign _GEN_788 = 5'h13 == _T_626_0 ? _GEN_7 : _T_18251_0_19;
  assign _GEN_789 = 5'h14 == _T_626_0 ? _GEN_7 : _T_18251_0_20;
  assign _GEN_790 = 5'h15 == _T_626_0 ? _GEN_7 : _T_18251_0_21;
  assign _GEN_791 = 5'h16 == _T_626_0 ? _GEN_7 : _T_18251_0_22;
  assign _GEN_792 = 5'h17 == _T_626_0 ? _GEN_7 : _T_18251_0_23;
  assign _GEN_793 = 5'h18 == _T_626_0 ? _GEN_7 : _T_18251_0_24;
  assign _GEN_794 = 5'h19 == _T_626_0 ? _GEN_7 : _T_18251_0_25;
  assign _GEN_795 = 5'h1a == _T_626_0 ? _GEN_7 : _T_18251_0_26;
  assign _GEN_796 = 5'h1b == _T_626_0 ? _GEN_7 : _T_18251_0_27;
  assign _GEN_797 = 5'h1c == _T_626_0 ? _GEN_7 : _T_18251_0_28;
  assign _GEN_798 = 5'h1d == _T_626_0 ? _GEN_7 : _T_18251_0_29;
  assign _GEN_799 = 5'h1e == _T_626_0 ? _GEN_7 : _T_18251_0_30;
  assign _GEN_800 = 5'h1f == _T_626_0 ? _GEN_7 : _T_18251_0_31;
  assign _GEN_801 = _T_614_0 ? _GEN_769 : _T_18251_0_0;
  assign _GEN_802 = _T_614_0 ? _GEN_770 : _T_18251_0_1;
  assign _GEN_803 = _T_614_0 ? _GEN_771 : _T_18251_0_2;
  assign _GEN_804 = _T_614_0 ? _GEN_772 : _T_18251_0_3;
  assign _GEN_805 = _T_614_0 ? _GEN_773 : _T_18251_0_4;
  assign _GEN_806 = _T_614_0 ? _GEN_774 : _T_18251_0_5;
  assign _GEN_807 = _T_614_0 ? _GEN_775 : _T_18251_0_6;
  assign _GEN_808 = _T_614_0 ? _GEN_776 : _T_18251_0_7;
  assign _GEN_809 = _T_614_0 ? _GEN_777 : _T_18251_0_8;
  assign _GEN_810 = _T_614_0 ? _GEN_778 : _T_18251_0_9;
  assign _GEN_811 = _T_614_0 ? _GEN_779 : _T_18251_0_10;
  assign _GEN_812 = _T_614_0 ? _GEN_780 : _T_18251_0_11;
  assign _GEN_813 = _T_614_0 ? _GEN_781 : _T_18251_0_12;
  assign _GEN_814 = _T_614_0 ? _GEN_782 : _T_18251_0_13;
  assign _GEN_815 = _T_614_0 ? _GEN_783 : _T_18251_0_14;
  assign _GEN_816 = _T_614_0 ? _GEN_784 : _T_18251_0_15;
  assign _GEN_817 = _T_614_0 ? _GEN_785 : _T_18251_0_16;
  assign _GEN_818 = _T_614_0 ? _GEN_786 : _T_18251_0_17;
  assign _GEN_819 = _T_614_0 ? _GEN_787 : _T_18251_0_18;
  assign _GEN_820 = _T_614_0 ? _GEN_788 : _T_18251_0_19;
  assign _GEN_821 = _T_614_0 ? _GEN_789 : _T_18251_0_20;
  assign _GEN_822 = _T_614_0 ? _GEN_790 : _T_18251_0_21;
  assign _GEN_823 = _T_614_0 ? _GEN_791 : _T_18251_0_22;
  assign _GEN_824 = _T_614_0 ? _GEN_792 : _T_18251_0_23;
  assign _GEN_825 = _T_614_0 ? _GEN_793 : _T_18251_0_24;
  assign _GEN_826 = _T_614_0 ? _GEN_794 : _T_18251_0_25;
  assign _GEN_827 = _T_614_0 ? _GEN_795 : _T_18251_0_26;
  assign _GEN_828 = _T_614_0 ? _GEN_796 : _T_18251_0_27;
  assign _GEN_829 = _T_614_0 ? _GEN_797 : _T_18251_0_28;
  assign _GEN_830 = _T_614_0 ? _GEN_798 : _T_18251_0_29;
  assign _GEN_831 = _T_614_0 ? _GEN_799 : _T_18251_0_30;
  assign _GEN_832 = _T_614_0 ? _GEN_800 : _T_18251_0_31;
  assign _T_18510 = _T_18494 & _T_608_0;
  assign _T_18513 = _T_18510 & _T_18170;
  assign _T_18519 = _T_18513 & _T_18496;
  assign _GEN_833 = _T_18519 ? 1'h1 : _T_18161_0;
  assign _GEN_834 = _T_18519 ? _T_602_0 : _T_18174_0;
  assign _T_18528 = _T_18483 == 1'h0;
  assign _T_18529 = _T_18161_0 & _T_18528;
  assign _T_18634 = {_T_18251_0_1,_T_18251_0_0};
  assign _T_18635 = {_T_18251_0_3,_T_18251_0_2};
  assign _T_18636 = {_T_18635,_T_18634};
  assign _T_18637 = {_T_18251_0_5,_T_18251_0_4};
  assign _T_18638 = {_T_18251_0_7,_T_18251_0_6};
  assign _T_18639 = {_T_18638,_T_18637};
  assign _T_18640 = {_T_18639,_T_18636};
  assign _T_18641 = {_T_18251_0_9,_T_18251_0_8};
  assign _T_18642 = {_T_18251_0_11,_T_18251_0_10};
  assign _T_18643 = {_T_18642,_T_18641};
  assign _T_18644 = {_T_18251_0_13,_T_18251_0_12};
  assign _T_18645 = {_T_18251_0_15,_T_18251_0_14};
  assign _T_18646 = {_T_18645,_T_18644};
  assign _T_18647 = {_T_18646,_T_18643};
  assign _T_18648 = {_T_18647,_T_18640};
  assign _T_18649 = {_T_18251_0_17,_T_18251_0_16};
  assign _T_18650 = {_T_18251_0_19,_T_18251_0_18};
  assign _T_18651 = {_T_18650,_T_18649};
  assign _T_18652 = {_T_18251_0_21,_T_18251_0_20};
  assign _T_18653 = {_T_18251_0_23,_T_18251_0_22};
  assign _T_18654 = {_T_18653,_T_18652};
  assign _T_18655 = {_T_18654,_T_18651};
  assign _T_18656 = {_T_18251_0_25,_T_18251_0_24};
  assign _T_18657 = {_T_18251_0_27,_T_18251_0_26};
  assign _T_18658 = {_T_18657,_T_18656};
  assign _T_18659 = {_T_18251_0_29,_T_18251_0_28};
  assign _T_18660 = {_T_18251_0_31,_T_18251_0_30};
  assign _T_18661 = {_T_18660,_T_18659};
  assign _T_18662 = {_T_18661,_T_18658};
  assign _T_18663 = {_T_18662,_T_18655};
  assign _T_18664 = {_T_18663,_T_18648};
  assign _T_18665 = _T_18664[511:0];
  assign _T_18668 = _T_18664[1023:512];
  assign _T_18669 = _T_18489 ? _T_18668 : _T_18665;
  assign _T_18676 = io_axi_outputMemAddrValids_3 & io_axi_outputMemAddrReadys_3;
  assign _T_18683 = _T_18492 & _T_18170;
  assign _T_18684 = _T_18676 | _T_18683;
  assign _T_18686 = _T_18480 == 1'h0;
  assign _T_18689 = _T_18480 + 1'h1;
  assign _T_18690 = _T_18689[0:0];
  assign _GEN_835 = _T_18686 ? 1'h1 : _T_18483;
  assign _GEN_836 = _T_18686 ? _T_18480 : _T_18690;
  assign _GEN_837 = _T_18684 ? _GEN_835 : _T_18483;
  assign _GEN_838 = _T_18684 ? _GEN_836 : _T_18480;
  assign _T_18691 = io_axi_outputMemBlockValids_3 & io_axi_outputMemBlockReadys_3;
  assign _T_18696 = _T_18489 + 1'h1;
  assign _T_18697 = _T_18696[0:0];
  assign _T_18698 = _T_18489 ? 1'h0 : _T_18697;
  assign _GEN_839 = _T_18691 ? _T_18698 : _T_18489;
  assign _T_18702 = _T_18691 & _T_18489;
  assign _T_18709 = _T_18486 < _T_18480;
  assign _T_18710 = _T_18709 | _T_18483;
  assign _T_18711 = _T_18170 & _T_18710;
  assign _T_18712 = _T_18702 | _T_18711;
  assign _T_18714 = _T_18486 == 1'h0;
  assign _T_18716 = _T_419 == 1'h0;
  assign _T_18719 = _T_419 + 1'h1;
  assign _T_18720 = _T_18719[0:0];
  assign _T_18721 = _T_18716 ? 1'h0 : _T_18720;
  assign _T_18730 = _T_18486 + 1'h1;
  assign _T_18731 = _T_18730[0:0];
  assign _GEN_840 = _T_18714 ? _T_18721 : _T_419;
  assign _GEN_841 = _T_18714 ? 1'h0 : _GEN_766;
  assign _GEN_842 = _T_18714 ? 1'h0 : _T_18731;
  assign _GEN_843 = _T_18714 ? 1'h0 : _GEN_838;
  assign _GEN_844 = _T_18714 ? 1'h0 : _GEN_837;
  assign _GEN_845 = _T_18714 ? 1'h0 : _GEN_767;
  assign _GEN_846 = _T_18714 ? 1'h0 : _GEN_833;
  assign _GEN_847 = _T_18714 ? 1'h0 : _GEN_768;
  assign _GEN_848 = _T_18712 ? _GEN_840 : _T_419;
  assign _GEN_849 = _T_18712 ? _GEN_841 : _GEN_766;
  assign _GEN_850 = _T_18712 ? _GEN_842 : _T_18486;
  assign _GEN_851 = _T_18712 ? _GEN_843 : _GEN_838;
  assign _GEN_852 = _T_18712 ? _GEN_844 : _GEN_837;
  assign _GEN_853 = _T_18712 ? _GEN_845 : _GEN_767;
  assign _GEN_854 = _T_18712 ? _GEN_846 : _GEN_833;
  assign _GEN_855 = _T_18712 ? _GEN_847 : _GEN_768;
  assign _T_18747 = _T_18716 ? _T_18519 : 1'h0;
  assign _T_18750 = _T_524_0 & _T_560_0;
  assign _T_18751 = _T_18750 & _T_596_0;
  assign _T_18752 = _T_18751 & _T_632_0;
  assign _T_18753 = _T_18752 & _T_16346;
  assign _T_18754 = _T_18753 & _T_16954;
  assign _T_18755 = _T_18754 & _T_17562;
  assign cumFinished = _T_18755 & _T_18170;
  assign io_axi_inputMemAddrs_0 = {{32'd0}, _T_422_0};
  assign io_axi_inputMemAddrs_1 = {{32'd0}, _T_440_0};
  assign io_axi_inputMemAddrs_2 = {{32'd0}, _T_458_0};
  assign io_axi_inputMemAddrs_3 = {{32'd0}, _T_476_0};
  assign io_axi_inputMemAddrValids_0 = _T_1033;
  assign io_axi_inputMemAddrValids_1 = _T_4953;
  assign io_axi_inputMemAddrValids_2 = _T_8873;
  assign io_axi_inputMemAddrValids_3 = _T_12793;
  assign io_axi_inputMemAddrLens_0 = 8'h1;
  assign io_axi_inputMemAddrLens_1 = 8'h1;
  assign io_axi_inputMemAddrLens_2 = 8'h1;
  assign io_axi_inputMemAddrLens_3 = 8'h1;
  assign io_axi_inputMemBlockReadys_0 = _T_4538;
  assign io_axi_inputMemBlockReadys_1 = _T_8458;
  assign io_axi_inputMemBlockReadys_2 = _T_12378;
  assign io_axi_inputMemBlockReadys_3 = _T_16298;
  assign io_axi_outputMemAddrs_0 = {{32'd0}, _T_16350_0};
  assign io_axi_outputMemAddrs_1 = {{32'd0}, _T_16958_0};
  assign io_axi_outputMemAddrs_2 = {{32'd0}, _T_17566_0};
  assign io_axi_outputMemAddrs_3 = {{32'd0}, _T_18174_0};
  assign io_axi_outputMemAddrValids_0 = _T_16705;
  assign io_axi_outputMemAddrValids_1 = _T_17313;
  assign io_axi_outputMemAddrValids_2 = _T_17921;
  assign io_axi_outputMemAddrValids_3 = _T_18529;
  assign io_axi_outputMemAddrLens_0 = 8'h1;
  assign io_axi_outputMemAddrLens_1 = 8'h1;
  assign io_axi_outputMemAddrLens_2 = 8'h1;
  assign io_axi_outputMemAddrLens_3 = 8'h1;
  assign io_axi_outputMemAddrIds_0 = {{15'd0}, _T_16656};
  assign io_axi_outputMemAddrIds_1 = {{15'd0}, _T_17264};
  assign io_axi_outputMemAddrIds_2 = {{15'd0}, _T_17872};
  assign io_axi_outputMemAddrIds_3 = {{15'd0}, _T_18480};
  assign io_axi_outputMemBlocks_0 = _T_16845;
  assign io_axi_outputMemBlocks_1 = _T_17453;
  assign io_axi_outputMemBlocks_2 = _T_18061;
  assign io_axi_outputMemBlocks_3 = _T_18669;
  assign io_axi_outputMemBlockValids_0 = _T_16646_0;
  assign io_axi_outputMemBlockValids_1 = _T_17254_0;
  assign io_axi_outputMemBlockValids_2 = _T_17862_0;
  assign io_axi_outputMemBlockValids_3 = _T_18470_0;
  assign io_axi_outputMemBlockLasts_0 = _T_16665;
  assign io_axi_outputMemBlockLasts_1 = _T_17273;
  assign io_axi_outputMemBlockLasts_2 = _T_17881;
  assign io_axi_outputMemBlockLasts_3 = _T_18489;
  assign io_axi_finished = cumFinished;
  assign io_streamingCores_0_metadataPtr = 32'h0;
  assign io_streamingCores_0_inputMemBlock = _GEN_0;
  assign io_streamingCores_0_inputMemIdx = _T_973_0;
  assign io_streamingCores_0_inputMemBlockValid = _T_4555;
  assign io_streamingCores_0_outputMemAddrReady = _T_16923;
  assign io_streamingCores_1_metadataPtr = 32'h0;
  assign io_streamingCores_1_inputMemBlock = _GEN_1;
  assign io_streamingCores_1_inputMemIdx = _T_4893_0;
  assign io_streamingCores_1_inputMemBlockValid = _T_8475;
  assign io_streamingCores_1_outputMemAddrReady = _T_17531;
  assign io_streamingCores_2_metadataPtr = 32'h0;
  assign io_streamingCores_2_inputMemBlock = _GEN_2;
  assign io_streamingCores_2_inputMemIdx = _T_8813_0;
  assign io_streamingCores_2_inputMemBlockValid = _T_12395;
  assign io_streamingCores_2_outputMemAddrReady = _T_18139;
  assign io_streamingCores_3_metadataPtr = 32'h0;
  assign io_streamingCores_3_inputMemBlock = _GEN_3;
  assign io_streamingCores_3_inputMemIdx = _T_12733_0;
  assign io_streamingCores_3_inputMemBlockValid = _T_16315;
  assign io_streamingCores_3_outputMemAddrReady = _T_18747;
  assign _T_422_0 = io_streamingCores_0_inputMemAddr;
  assign _T_428_0 = io_streamingCores_0_inputMemAddrValid;
  assign _T_434_0 = io_streamingCores_0_inputMemAddrsFinished;
  assign _T_440_0 = io_streamingCores_1_inputMemAddr;
  assign _T_446_0 = io_streamingCores_1_inputMemAddrValid;
  assign _T_452_0 = io_streamingCores_1_inputMemAddrsFinished;
  assign _T_458_0 = io_streamingCores_2_inputMemAddr;
  assign _T_464_0 = io_streamingCores_2_inputMemAddrValid;
  assign _T_470_0 = io_streamingCores_2_inputMemAddrsFinished;
  assign _T_476_0 = io_streamingCores_3_inputMemAddr;
  assign _T_482_0 = io_streamingCores_3_inputMemAddrValid;
  assign _T_488_0 = io_streamingCores_3_inputMemAddrsFinished;
  assign _T_494_0 = io_streamingCores_0_outputMemAddr;
  assign _T_500_0 = io_streamingCores_0_outputMemAddrValid;
  assign _T_506_0 = io_streamingCores_0_outputMemBlockValid;
  assign _T_512_0 = io_streamingCores_0_outputMemBlock;
  assign _T_518_0 = io_streamingCores_0_outputMemIdx;
  assign _T_524_0 = io_streamingCores_0_outputFinished;
  assign _T_530_0 = io_streamingCores_1_outputMemAddr;
  assign _T_536_0 = io_streamingCores_1_outputMemAddrValid;
  assign _T_542_0 = io_streamingCores_1_outputMemBlockValid;
  assign _T_548_0 = io_streamingCores_1_outputMemBlock;
  assign _T_554_0 = io_streamingCores_1_outputMemIdx;
  assign _T_560_0 = io_streamingCores_1_outputFinished;
  assign _T_566_0 = io_streamingCores_2_outputMemAddr;
  assign _T_572_0 = io_streamingCores_2_outputMemAddrValid;
  assign _T_578_0 = io_streamingCores_2_outputMemBlockValid;
  assign _T_584_0 = io_streamingCores_2_outputMemBlock;
  assign _T_590_0 = io_streamingCores_2_outputMemIdx;
  assign _T_596_0 = io_streamingCores_2_outputFinished;
  assign _T_602_0 = io_streamingCores_3_outputMemAddr;
  assign _T_608_0 = io_streamingCores_3_outputMemAddrValid;
  assign _T_614_0 = io_streamingCores_3_outputMemBlockValid;
  assign _T_620_0 = io_streamingCores_3_outputMemBlock;
  assign _T_626_0 = io_streamingCores_3_outputMemIdx;
  assign _T_632_0 = io_streamingCores_3_outputFinished;
  assign _GEN_0 = _GEN_129;
  assign _GEN_1 = _GEN_251;
  assign _GEN_2 = _GEN_373;
  assign _GEN_3 = _GEN_495;
  assign _GEN_4 = _T_512_0;
  assign _GEN_5 = _T_548_0;
  assign _GEN_6 = _T_584_0;
  assign _GEN_7 = _T_620_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_389 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_395 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_401 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_407 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_410 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_413 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_416 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_419 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_638 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_652_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_673_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_754_0_0 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_754_0_1 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_754_0_2 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_754_0_3 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_754_0_4 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_754_0_5 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_754_0_6 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_754_0_7 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_754_0_8 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_754_0_9 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_754_0_10 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_754_0_11 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_754_0_12 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_754_0_13 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_754_0_14 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_754_0_15 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_754_0_16 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_754_0_17 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_754_0_18 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_754_0_19 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_754_0_20 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_754_0_21 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_754_0_22 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_754_0_23 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_754_0_24 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_754_0_25 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_754_0_26 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_754_0_27 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_754_0_28 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_754_0_29 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_754_0_30 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_754_0_31 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_973_0 = _RAND_43[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_994_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_1004 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_1007 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_1010 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_4558 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_4572_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_4593_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_4674_0_0 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_4674_0_1 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_4674_0_2 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_4674_0_3 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_4674_0_4 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_4674_0_5 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_4674_0_6 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_4674_0_7 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_4674_0_8 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_4674_0_9 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_4674_0_10 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_4674_0_11 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_4674_0_12 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_4674_0_13 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_4674_0_14 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_4674_0_15 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_4674_0_16 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_4674_0_17 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_4674_0_18 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_4674_0_19 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_4674_0_20 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_4674_0_21 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_4674_0_22 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_4674_0_23 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_4674_0_24 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_4674_0_25 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_4674_0_26 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_4674_0_27 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_4674_0_28 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_4674_0_29 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_4674_0_30 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_4674_0_31 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_4893_0 = _RAND_83[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_4914_0 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_4924 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_4927 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_4930 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_8478 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_8492_0 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_8513_0 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_8594_0_0 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_8594_0_1 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_8594_0_2 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_8594_0_3 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_8594_0_4 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_8594_0_5 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_8594_0_6 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_8594_0_7 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_8594_0_8 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_8594_0_9 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_8594_0_10 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_8594_0_11 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_8594_0_12 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_8594_0_13 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_8594_0_14 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_8594_0_15 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_8594_0_16 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_8594_0_17 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_8594_0_18 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_8594_0_19 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_8594_0_20 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_8594_0_21 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_8594_0_22 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_8594_0_23 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_8594_0_24 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_8594_0_25 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_8594_0_26 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_8594_0_27 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_8594_0_28 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_8594_0_29 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_8594_0_30 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_8594_0_31 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_8813_0 = _RAND_123[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_8834_0 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_8844 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_8847 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_8850 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_12398 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_12412_0 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_12433_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_12514_0_0 = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_12514_0_1 = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_12514_0_2 = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_12514_0_3 = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  _T_12514_0_4 = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_12514_0_5 = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  _T_12514_0_6 = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  _T_12514_0_7 = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  _T_12514_0_8 = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  _T_12514_0_9 = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  _T_12514_0_10 = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  _T_12514_0_11 = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  _T_12514_0_12 = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  _T_12514_0_13 = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  _T_12514_0_14 = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  _T_12514_0_15 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  _T_12514_0_16 = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  _T_12514_0_17 = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  _T_12514_0_18 = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  _T_12514_0_19 = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  _T_12514_0_20 = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  _T_12514_0_21 = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  _T_12514_0_22 = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  _T_12514_0_23 = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _T_12514_0_24 = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  _T_12514_0_25 = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _T_12514_0_26 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  _T_12514_0_27 = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  _T_12514_0_28 = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _T_12514_0_29 = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  _T_12514_0_30 = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  _T_12514_0_31 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  _T_12733_0 = _RAND_163[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  _T_12754_0 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  _T_12764 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  _T_12767 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  _T_12770 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  _T_16318 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  _T_16337_0 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  _T_16350_0 = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  _T_16427_0_0 = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  _T_16427_0_1 = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  _T_16427_0_2 = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  _T_16427_0_3 = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  _T_16427_0_4 = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  _T_16427_0_5 = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  _T_16427_0_6 = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  _T_16427_0_7 = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  _T_16427_0_8 = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  _T_16427_0_9 = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  _T_16427_0_10 = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  _T_16427_0_11 = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  _T_16427_0_12 = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  _T_16427_0_13 = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  _T_16427_0_14 = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  _T_16427_0_15 = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  _T_16427_0_16 = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  _T_16427_0_17 = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  _T_16427_0_18 = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  _T_16427_0_19 = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  _T_16427_0_20 = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  _T_16427_0_21 = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  _T_16427_0_22 = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  _T_16427_0_23 = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  _T_16427_0_24 = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  _T_16427_0_25 = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  _T_16427_0_26 = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  _T_16427_0_27 = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  _T_16427_0_28 = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  _T_16427_0_29 = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  _T_16427_0_30 = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  _T_16427_0_31 = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  _T_16646_0 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  _T_16656 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  _T_16659 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  _T_16662 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  _T_16665 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  _T_16668 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  _T_16926 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  _T_16945_0 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  _T_16958_0 = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  _T_17035_0_0 = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  _T_17035_0_1 = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  _T_17035_0_2 = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  _T_17035_0_3 = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  _T_17035_0_4 = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  _T_17035_0_5 = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  _T_17035_0_6 = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  _T_17035_0_7 = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  _T_17035_0_8 = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  _T_17035_0_9 = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  _T_17035_0_10 = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  _T_17035_0_11 = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  _T_17035_0_12 = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  _T_17035_0_13 = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  _T_17035_0_14 = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  _T_17035_0_15 = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  _T_17035_0_16 = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  _T_17035_0_17 = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  _T_17035_0_18 = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  _T_17035_0_19 = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  _T_17035_0_20 = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  _T_17035_0_21 = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  _T_17035_0_22 = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  _T_17035_0_23 = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  _T_17035_0_24 = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  _T_17035_0_25 = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  _T_17035_0_26 = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  _T_17035_0_27 = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  _T_17035_0_28 = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  _T_17035_0_29 = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  _T_17035_0_30 = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  _T_17035_0_31 = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  _T_17254_0 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  _T_17264 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  _T_17267 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  _T_17270 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  _T_17273 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{$random}};
  _T_17276 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{$random}};
  _T_17534 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{$random}};
  _T_17553_0 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{$random}};
  _T_17566_0 = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{$random}};
  _T_17643_0_0 = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{$random}};
  _T_17643_0_1 = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{$random}};
  _T_17643_0_2 = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{$random}};
  _T_17643_0_3 = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{$random}};
  _T_17643_0_4 = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{$random}};
  _T_17643_0_5 = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{$random}};
  _T_17643_0_6 = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{$random}};
  _T_17643_0_7 = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{$random}};
  _T_17643_0_8 = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{$random}};
  _T_17643_0_9 = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{$random}};
  _T_17643_0_10 = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{$random}};
  _T_17643_0_11 = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{$random}};
  _T_17643_0_12 = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{$random}};
  _T_17643_0_13 = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{$random}};
  _T_17643_0_14 = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{$random}};
  _T_17643_0_15 = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{$random}};
  _T_17643_0_16 = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{$random}};
  _T_17643_0_17 = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{$random}};
  _T_17643_0_18 = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{$random}};
  _T_17643_0_19 = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{$random}};
  _T_17643_0_20 = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{$random}};
  _T_17643_0_21 = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{$random}};
  _T_17643_0_22 = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{$random}};
  _T_17643_0_23 = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{$random}};
  _T_17643_0_24 = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{$random}};
  _T_17643_0_25 = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{$random}};
  _T_17643_0_26 = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{$random}};
  _T_17643_0_27 = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{$random}};
  _T_17643_0_28 = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{$random}};
  _T_17643_0_29 = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{$random}};
  _T_17643_0_30 = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{$random}};
  _T_17643_0_31 = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{$random}};
  _T_17862_0 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{$random}};
  _T_17872 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{$random}};
  _T_17875 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{$random}};
  _T_17878 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{$random}};
  _T_17881 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{$random}};
  _T_17884 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{$random}};
  _T_18142 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{$random}};
  _T_18161_0 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{$random}};
  _T_18174_0 = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{$random}};
  _T_18251_0_0 = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{$random}};
  _T_18251_0_1 = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{$random}};
  _T_18251_0_2 = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{$random}};
  _T_18251_0_3 = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{$random}};
  _T_18251_0_4 = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{$random}};
  _T_18251_0_5 = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{$random}};
  _T_18251_0_6 = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{$random}};
  _T_18251_0_7 = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{$random}};
  _T_18251_0_8 = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{$random}};
  _T_18251_0_9 = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{$random}};
  _T_18251_0_10 = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{$random}};
  _T_18251_0_11 = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{$random}};
  _T_18251_0_12 = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{$random}};
  _T_18251_0_13 = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{$random}};
  _T_18251_0_14 = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{$random}};
  _T_18251_0_15 = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{$random}};
  _T_18251_0_16 = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{$random}};
  _T_18251_0_17 = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{$random}};
  _T_18251_0_18 = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{$random}};
  _T_18251_0_19 = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{$random}};
  _T_18251_0_20 = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{$random}};
  _T_18251_0_21 = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{$random}};
  _T_18251_0_22 = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{$random}};
  _T_18251_0_23 = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{$random}};
  _T_18251_0_24 = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{$random}};
  _T_18251_0_25 = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{$random}};
  _T_18251_0_26 = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{$random}};
  _T_18251_0_27 = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{$random}};
  _T_18251_0_28 = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{$random}};
  _T_18251_0_29 = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{$random}};
  _T_18251_0_30 = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{$random}};
  _T_18251_0_31 = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{$random}};
  _T_18470_0 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{$random}};
  _T_18480 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{$random}};
  _T_18483 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{$random}};
  _T_18486 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{$random}};
  _T_18489 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{$random}};
  _T_18492 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_389 <= 1'h0;
    end else begin
      if (_T_4504) begin
        if (_T_4516) begin
          if (_T_4518) begin
            _T_389 <= 1'h0;
          end else begin
            _T_389 <= _T_4522;
          end
        end
      end
    end
    if (reset) begin
      _T_395 <= 1'h0;
    end else begin
      if (_T_8424) begin
        if (_T_8436) begin
          if (_T_8438) begin
            _T_395 <= 1'h0;
          end else begin
            _T_395 <= _T_8442;
          end
        end
      end
    end
    if (reset) begin
      _T_401 <= 1'h0;
    end else begin
      if (_T_12344) begin
        if (_T_12356) begin
          if (_T_12358) begin
            _T_401 <= 1'h0;
          end else begin
            _T_401 <= _T_12362;
          end
        end
      end
    end
    if (reset) begin
      _T_407 <= 1'h0;
    end else begin
      if (_T_16264) begin
        if (_T_16276) begin
          if (_T_16278) begin
            _T_407 <= 1'h0;
          end else begin
            _T_407 <= _T_16282;
          end
        end
      end
    end
    if (reset) begin
      _T_410 <= 1'h0;
    end else begin
      if (_T_16888) begin
        if (_T_16890) begin
          if (_T_16892) begin
            _T_410 <= 1'h0;
          end else begin
            _T_410 <= _T_16896;
          end
        end
      end
    end
    if (reset) begin
      _T_413 <= 1'h0;
    end else begin
      if (_T_17496) begin
        if (_T_17498) begin
          if (_T_17500) begin
            _T_413 <= 1'h0;
          end else begin
            _T_413 <= _T_17504;
          end
        end
      end
    end
    if (reset) begin
      _T_416 <= 1'h0;
    end else begin
      if (_T_18104) begin
        if (_T_18106) begin
          if (_T_18108) begin
            _T_416 <= 1'h0;
          end else begin
            _T_416 <= _T_18112;
          end
        end
      end
    end
    if (reset) begin
      _T_419 <= 1'h0;
    end else begin
      if (_T_18712) begin
        if (_T_18714) begin
          if (_T_18716) begin
            _T_419 <= 1'h0;
          end else begin
            _T_419 <= _T_18720;
          end
        end
      end
    end
    if (reset) begin
      _T_638 <= 1'h0;
    end else begin
      if (_T_1048) begin
        if (_T_1060) begin
          _T_638 <= 1'h0;
        end else begin
          if (_T_1016) begin
            _T_638 <= _T_1019;
          end
        end
      end else begin
        if (_T_1016) begin
          _T_638 <= _T_1019;
        end
      end
    end
    if (reset) begin
      _T_652_0 <= 1'h0;
    end else begin
      if (_T_4504) begin
        if (io_axi_inputMemBlockReadys_0) begin
          if (_T_994_0) begin
            if (_T_1074) begin
              _T_652_0 <= 1'h0;
            end else begin
              if (_T_1048) begin
                _T_652_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_1048) begin
              _T_652_0 <= 1'h1;
            end
          end
        end else begin
          _T_652_0 <= 1'h0;
        end
      end else begin
        if (_T_994_0) begin
          if (_T_1074) begin
            _T_652_0 <= 1'h0;
          end else begin
            if (_T_1048) begin
              _T_652_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_1048) begin
            _T_652_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_673_0 <= 1'h0;
    end else begin
      if (_T_994_0) begin
        if (_T_1074) begin
          _T_673_0 <= 1'h0;
        end else begin
          if (_T_1048) begin
            if (io_axi_inputMemAddrValids_0) begin
              _T_673_0 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_1048) begin
          if (io_axi_inputMemAddrValids_0) begin
            _T_673_0 <= 1'h1;
          end
        end
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_0 <= _T_1195;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_1 <= _T_1301;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_2 <= _T_1407;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_3 <= _T_1513;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_4 <= _T_1619;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_5 <= _T_1725;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_6 <= _T_1831;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_7 <= _T_1937;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_8 <= _T_2043;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_9 <= _T_2149;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_10 <= _T_2255;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_11 <= _T_2361;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_12 <= _T_2467;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_13 <= _T_2573;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_14 <= _T_2679;
      end
    end
    if (_T_1082) begin
      if (_T_1091) begin
        _T_754_0_15 <= _T_2785;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_16 <= _T_1195;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_17 <= _T_1301;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_18 <= _T_1407;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_19 <= _T_1513;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_20 <= _T_1619;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_21 <= _T_1725;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_22 <= _T_1831;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_23 <= _T_1937;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_24 <= _T_2043;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_25 <= _T_2149;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_26 <= _T_2255;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_27 <= _T_2361;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_28 <= _T_2467;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_29 <= _T_2573;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_30 <= _T_2679;
      end
    end
    if (_T_1082) begin
      if (_T_1010) begin
        _T_754_0_31 <= _T_2785;
      end
    end
    if (reset) begin
      _T_973_0 <= 5'h0;
    end else begin
      if (_T_994_0) begin
        if (_T_1074) begin
          _T_973_0 <= 5'h0;
        end else begin
          _T_973_0 <= _T_1081;
        end
      end
    end
    if (reset) begin
      _T_994_0 <= 1'h0;
    end else begin
      if (_T_4504) begin
        if (io_axi_inputMemBlockReadys_0) begin
          _T_994_0 <= 1'h1;
        end else begin
          if (_T_994_0) begin
            if (_T_1074) begin
              _T_994_0 <= 1'h0;
            end
          end
        end
      end else begin
        if (_T_994_0) begin
          if (_T_1074) begin
            _T_994_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_1004 <= 1'h0;
    end else begin
      if (_T_1048) begin
        if (_T_1060) begin
          _T_1004 <= 1'h0;
        end else begin
          _T_1004 <= _T_1072;
        end
      end
    end
    if (reset) begin
      _T_1007 <= 1'h0;
    end else begin
      if (_T_4504) begin
        if (_T_4516) begin
          _T_1007 <= 1'h0;
        end else begin
          _T_1007 <= _T_4527;
        end
      end
    end
    if (reset) begin
      _T_1010 <= 1'h0;
    end else begin
      if (_T_1082) begin
        if (_T_1010) begin
          _T_1010 <= 1'h0;
        end else begin
          _T_1010 <= _T_1088;
        end
      end
    end
    if (reset) begin
      _T_4558 <= 1'h0;
    end else begin
      if (_T_4968) begin
        if (_T_4980) begin
          _T_4558 <= 1'h0;
        end else begin
          if (_T_4936) begin
            _T_4558 <= _T_4939;
          end
        end
      end else begin
        if (_T_4936) begin
          _T_4558 <= _T_4939;
        end
      end
    end
    if (reset) begin
      _T_4572_0 <= 1'h0;
    end else begin
      if (_T_8424) begin
        if (io_axi_inputMemBlockReadys_1) begin
          if (_T_4914_0) begin
            if (_T_4994) begin
              _T_4572_0 <= 1'h0;
            end else begin
              if (_T_4968) begin
                _T_4572_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_4968) begin
              _T_4572_0 <= 1'h1;
            end
          end
        end else begin
          _T_4572_0 <= 1'h0;
        end
      end else begin
        if (_T_4914_0) begin
          if (_T_4994) begin
            _T_4572_0 <= 1'h0;
          end else begin
            if (_T_4968) begin
              _T_4572_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_4968) begin
            _T_4572_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_4593_0 <= 1'h0;
    end else begin
      if (_T_4914_0) begin
        if (_T_4994) begin
          _T_4593_0 <= 1'h0;
        end else begin
          if (_T_4968) begin
            if (io_axi_inputMemAddrValids_1) begin
              _T_4593_0 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_4968) begin
          if (io_axi_inputMemAddrValids_1) begin
            _T_4593_0 <= 1'h1;
          end
        end
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_0 <= _T_5115;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_1 <= _T_5221;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_2 <= _T_5327;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_3 <= _T_5433;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_4 <= _T_5539;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_5 <= _T_5645;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_6 <= _T_5751;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_7 <= _T_5857;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_8 <= _T_5963;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_9 <= _T_6069;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_10 <= _T_6175;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_11 <= _T_6281;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_12 <= _T_6387;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_13 <= _T_6493;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_14 <= _T_6599;
      end
    end
    if (_T_5002) begin
      if (_T_5011) begin
        _T_4674_0_15 <= _T_6705;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_16 <= _T_5115;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_17 <= _T_5221;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_18 <= _T_5327;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_19 <= _T_5433;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_20 <= _T_5539;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_21 <= _T_5645;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_22 <= _T_5751;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_23 <= _T_5857;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_24 <= _T_5963;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_25 <= _T_6069;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_26 <= _T_6175;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_27 <= _T_6281;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_28 <= _T_6387;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_29 <= _T_6493;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_30 <= _T_6599;
      end
    end
    if (_T_5002) begin
      if (_T_4930) begin
        _T_4674_0_31 <= _T_6705;
      end
    end
    if (reset) begin
      _T_4893_0 <= 5'h0;
    end else begin
      if (_T_4914_0) begin
        if (_T_4994) begin
          _T_4893_0 <= 5'h0;
        end else begin
          _T_4893_0 <= _T_5001;
        end
      end
    end
    if (reset) begin
      _T_4914_0 <= 1'h0;
    end else begin
      if (_T_8424) begin
        if (io_axi_inputMemBlockReadys_1) begin
          _T_4914_0 <= 1'h1;
        end else begin
          if (_T_4914_0) begin
            if (_T_4994) begin
              _T_4914_0 <= 1'h0;
            end
          end
        end
      end else begin
        if (_T_4914_0) begin
          if (_T_4994) begin
            _T_4914_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_4924 <= 1'h0;
    end else begin
      if (_T_4968) begin
        if (_T_4980) begin
          _T_4924 <= 1'h0;
        end else begin
          _T_4924 <= _T_4992;
        end
      end
    end
    if (reset) begin
      _T_4927 <= 1'h0;
    end else begin
      if (_T_8424) begin
        if (_T_8436) begin
          _T_4927 <= 1'h0;
        end else begin
          _T_4927 <= _T_8447;
        end
      end
    end
    if (reset) begin
      _T_4930 <= 1'h0;
    end else begin
      if (_T_5002) begin
        if (_T_4930) begin
          _T_4930 <= 1'h0;
        end else begin
          _T_4930 <= _T_5008;
        end
      end
    end
    if (reset) begin
      _T_8478 <= 1'h0;
    end else begin
      if (_T_8888) begin
        if (_T_8900) begin
          _T_8478 <= 1'h0;
        end else begin
          if (_T_8856) begin
            _T_8478 <= _T_8859;
          end
        end
      end else begin
        if (_T_8856) begin
          _T_8478 <= _T_8859;
        end
      end
    end
    if (reset) begin
      _T_8492_0 <= 1'h0;
    end else begin
      if (_T_12344) begin
        if (io_axi_inputMemBlockReadys_2) begin
          if (_T_8834_0) begin
            if (_T_8914) begin
              _T_8492_0 <= 1'h0;
            end else begin
              if (_T_8888) begin
                _T_8492_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_8888) begin
              _T_8492_0 <= 1'h1;
            end
          end
        end else begin
          _T_8492_0 <= 1'h0;
        end
      end else begin
        if (_T_8834_0) begin
          if (_T_8914) begin
            _T_8492_0 <= 1'h0;
          end else begin
            if (_T_8888) begin
              _T_8492_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_8888) begin
            _T_8492_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_8513_0 <= 1'h0;
    end else begin
      if (_T_8834_0) begin
        if (_T_8914) begin
          _T_8513_0 <= 1'h0;
        end else begin
          if (_T_8888) begin
            if (io_axi_inputMemAddrValids_2) begin
              _T_8513_0 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_8888) begin
          if (io_axi_inputMemAddrValids_2) begin
            _T_8513_0 <= 1'h1;
          end
        end
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_0 <= _T_9035;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_1 <= _T_9141;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_2 <= _T_9247;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_3 <= _T_9353;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_4 <= _T_9459;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_5 <= _T_9565;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_6 <= _T_9671;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_7 <= _T_9777;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_8 <= _T_9883;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_9 <= _T_9989;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_10 <= _T_10095;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_11 <= _T_10201;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_12 <= _T_10307;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_13 <= _T_10413;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_14 <= _T_10519;
      end
    end
    if (_T_8922) begin
      if (_T_8931) begin
        _T_8594_0_15 <= _T_10625;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_16 <= _T_9035;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_17 <= _T_9141;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_18 <= _T_9247;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_19 <= _T_9353;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_20 <= _T_9459;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_21 <= _T_9565;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_22 <= _T_9671;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_23 <= _T_9777;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_24 <= _T_9883;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_25 <= _T_9989;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_26 <= _T_10095;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_27 <= _T_10201;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_28 <= _T_10307;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_29 <= _T_10413;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_30 <= _T_10519;
      end
    end
    if (_T_8922) begin
      if (_T_8850) begin
        _T_8594_0_31 <= _T_10625;
      end
    end
    if (reset) begin
      _T_8813_0 <= 5'h0;
    end else begin
      if (_T_8834_0) begin
        if (_T_8914) begin
          _T_8813_0 <= 5'h0;
        end else begin
          _T_8813_0 <= _T_8921;
        end
      end
    end
    if (reset) begin
      _T_8834_0 <= 1'h0;
    end else begin
      if (_T_12344) begin
        if (io_axi_inputMemBlockReadys_2) begin
          _T_8834_0 <= 1'h1;
        end else begin
          if (_T_8834_0) begin
            if (_T_8914) begin
              _T_8834_0 <= 1'h0;
            end
          end
        end
      end else begin
        if (_T_8834_0) begin
          if (_T_8914) begin
            _T_8834_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_8844 <= 1'h0;
    end else begin
      if (_T_8888) begin
        if (_T_8900) begin
          _T_8844 <= 1'h0;
        end else begin
          _T_8844 <= _T_8912;
        end
      end
    end
    if (reset) begin
      _T_8847 <= 1'h0;
    end else begin
      if (_T_12344) begin
        if (_T_12356) begin
          _T_8847 <= 1'h0;
        end else begin
          _T_8847 <= _T_12367;
        end
      end
    end
    if (reset) begin
      _T_8850 <= 1'h0;
    end else begin
      if (_T_8922) begin
        if (_T_8850) begin
          _T_8850 <= 1'h0;
        end else begin
          _T_8850 <= _T_8928;
        end
      end
    end
    if (reset) begin
      _T_12398 <= 1'h0;
    end else begin
      if (_T_12808) begin
        if (_T_12820) begin
          _T_12398 <= 1'h0;
        end else begin
          if (_T_12776) begin
            _T_12398 <= _T_12779;
          end
        end
      end else begin
        if (_T_12776) begin
          _T_12398 <= _T_12779;
        end
      end
    end
    if (reset) begin
      _T_12412_0 <= 1'h0;
    end else begin
      if (_T_16264) begin
        if (io_axi_inputMemBlockReadys_3) begin
          if (_T_12754_0) begin
            if (_T_12834) begin
              _T_12412_0 <= 1'h0;
            end else begin
              if (_T_12808) begin
                _T_12412_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_12808) begin
              _T_12412_0 <= 1'h1;
            end
          end
        end else begin
          _T_12412_0 <= 1'h0;
        end
      end else begin
        if (_T_12754_0) begin
          if (_T_12834) begin
            _T_12412_0 <= 1'h0;
          end else begin
            if (_T_12808) begin
              _T_12412_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_12808) begin
            _T_12412_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_12433_0 <= 1'h0;
    end else begin
      if (_T_12754_0) begin
        if (_T_12834) begin
          _T_12433_0 <= 1'h0;
        end else begin
          if (_T_12808) begin
            if (io_axi_inputMemAddrValids_3) begin
              _T_12433_0 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_12808) begin
          if (io_axi_inputMemAddrValids_3) begin
            _T_12433_0 <= 1'h1;
          end
        end
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_0 <= _T_12955;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_1 <= _T_13061;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_2 <= _T_13167;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_3 <= _T_13273;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_4 <= _T_13379;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_5 <= _T_13485;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_6 <= _T_13591;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_7 <= _T_13697;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_8 <= _T_13803;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_9 <= _T_13909;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_10 <= _T_14015;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_11 <= _T_14121;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_12 <= _T_14227;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_13 <= _T_14333;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_14 <= _T_14439;
      end
    end
    if (_T_12842) begin
      if (_T_12851) begin
        _T_12514_0_15 <= _T_14545;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_16 <= _T_12955;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_17 <= _T_13061;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_18 <= _T_13167;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_19 <= _T_13273;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_20 <= _T_13379;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_21 <= _T_13485;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_22 <= _T_13591;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_23 <= _T_13697;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_24 <= _T_13803;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_25 <= _T_13909;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_26 <= _T_14015;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_27 <= _T_14121;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_28 <= _T_14227;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_29 <= _T_14333;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_30 <= _T_14439;
      end
    end
    if (_T_12842) begin
      if (_T_12770) begin
        _T_12514_0_31 <= _T_14545;
      end
    end
    if (reset) begin
      _T_12733_0 <= 5'h0;
    end else begin
      if (_T_12754_0) begin
        if (_T_12834) begin
          _T_12733_0 <= 5'h0;
        end else begin
          _T_12733_0 <= _T_12841;
        end
      end
    end
    if (reset) begin
      _T_12754_0 <= 1'h0;
    end else begin
      if (_T_16264) begin
        if (io_axi_inputMemBlockReadys_3) begin
          _T_12754_0 <= 1'h1;
        end else begin
          if (_T_12754_0) begin
            if (_T_12834) begin
              _T_12754_0 <= 1'h0;
            end
          end
        end
      end else begin
        if (_T_12754_0) begin
          if (_T_12834) begin
            _T_12754_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_12764 <= 1'h0;
    end else begin
      if (_T_12808) begin
        if (_T_12820) begin
          _T_12764 <= 1'h0;
        end else begin
          _T_12764 <= _T_12832;
        end
      end
    end
    if (reset) begin
      _T_12767 <= 1'h0;
    end else begin
      if (_T_16264) begin
        if (_T_16276) begin
          _T_12767 <= 1'h0;
        end else begin
          _T_12767 <= _T_16287;
        end
      end
    end
    if (reset) begin
      _T_12770 <= 1'h0;
    end else begin
      if (_T_12842) begin
        if (_T_12770) begin
          _T_12770 <= 1'h0;
        end else begin
          _T_12770 <= _T_12848;
        end
      end
    end
    if (reset) begin
      _T_16318 <= 1'h0;
    end else begin
      if (_T_16888) begin
        if (_T_16890) begin
          _T_16318 <= 1'h0;
        end else begin
          if (_T_16318) begin
            _T_16318 <= _T_16323;
          end
        end
      end else begin
        if (_T_16318) begin
          _T_16318 <= _T_16323;
        end
      end
    end
    if (reset) begin
      _T_16337_0 <= 1'h0;
    end else begin
      if (_T_16888) begin
        if (_T_16890) begin
          _T_16337_0 <= 1'h0;
        end else begin
          if (_T_16695) begin
            _T_16337_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_16695) begin
          _T_16337_0 <= 1'h1;
        end
      end
    end
    if (_T_16695) begin
      _T_16350_0 <= _T_494_0;
    end
    if (_T_506_0) begin
      if (5'h0 == _T_518_0) begin
        _T_16427_0_0 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h1 == _T_518_0) begin
        _T_16427_0_1 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h2 == _T_518_0) begin
        _T_16427_0_2 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h3 == _T_518_0) begin
        _T_16427_0_3 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h4 == _T_518_0) begin
        _T_16427_0_4 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h5 == _T_518_0) begin
        _T_16427_0_5 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h6 == _T_518_0) begin
        _T_16427_0_6 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h7 == _T_518_0) begin
        _T_16427_0_7 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h8 == _T_518_0) begin
        _T_16427_0_8 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h9 == _T_518_0) begin
        _T_16427_0_9 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'ha == _T_518_0) begin
        _T_16427_0_10 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'hb == _T_518_0) begin
        _T_16427_0_11 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'hc == _T_518_0) begin
        _T_16427_0_12 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'hd == _T_518_0) begin
        _T_16427_0_13 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'he == _T_518_0) begin
        _T_16427_0_14 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'hf == _T_518_0) begin
        _T_16427_0_15 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h10 == _T_518_0) begin
        _T_16427_0_16 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h11 == _T_518_0) begin
        _T_16427_0_17 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h12 == _T_518_0) begin
        _T_16427_0_18 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h13 == _T_518_0) begin
        _T_16427_0_19 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h14 == _T_518_0) begin
        _T_16427_0_20 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h15 == _T_518_0) begin
        _T_16427_0_21 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h16 == _T_518_0) begin
        _T_16427_0_22 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h17 == _T_518_0) begin
        _T_16427_0_23 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h18 == _T_518_0) begin
        _T_16427_0_24 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h19 == _T_518_0) begin
        _T_16427_0_25 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h1a == _T_518_0) begin
        _T_16427_0_26 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h1b == _T_518_0) begin
        _T_16427_0_27 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h1c == _T_518_0) begin
        _T_16427_0_28 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h1d == _T_518_0) begin
        _T_16427_0_29 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h1e == _T_518_0) begin
        _T_16427_0_30 <= _GEN_4;
      end
    end
    if (_T_506_0) begin
      if (5'h1f == _T_518_0) begin
        _T_16427_0_31 <= _GEN_4;
      end
    end
    if (reset) begin
      _T_16646_0 <= 1'h0;
    end else begin
      if (_T_16888) begin
        if (_T_16890) begin
          _T_16646_0 <= 1'h0;
        end else begin
          if (_T_16680) begin
            _T_16646_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_16680) begin
          _T_16646_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_16656 <= 1'h0;
    end else begin
      if (_T_16888) begin
        if (_T_16890) begin
          _T_16656 <= 1'h0;
        end else begin
          if (_T_16860) begin
            if (!(_T_16862)) begin
              _T_16656 <= _T_16866;
            end
          end
        end
      end else begin
        if (_T_16860) begin
          if (!(_T_16862)) begin
            _T_16656 <= _T_16866;
          end
        end
      end
    end
    if (reset) begin
      _T_16659 <= 1'h0;
    end else begin
      if (_T_16888) begin
        if (_T_16890) begin
          _T_16659 <= 1'h0;
        end else begin
          if (_T_16860) begin
            if (_T_16862) begin
              _T_16659 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_16860) begin
          if (_T_16862) begin
            _T_16659 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_16662 <= 1'h0;
    end else begin
      if (_T_16888) begin
        if (_T_16890) begin
          _T_16662 <= 1'h0;
        end else begin
          _T_16662 <= _T_16907;
        end
      end
    end
    if (reset) begin
      _T_16665 <= 1'h0;
    end else begin
      if (_T_16867) begin
        if (_T_16665) begin
          _T_16665 <= 1'h0;
        end else begin
          _T_16665 <= _T_16873;
        end
      end
    end
    if (reset) begin
      _T_16668 <= 1'h0;
    end else begin
      if (_T_16888) begin
        if (_T_16890) begin
          _T_16668 <= 1'h0;
        end else begin
          if (_T_16673) begin
            _T_16668 <= 1'h1;
          end
        end
      end else begin
        if (_T_16673) begin
          _T_16668 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_16926 <= 1'h0;
    end else begin
      if (_T_17496) begin
        if (_T_17498) begin
          _T_16926 <= 1'h0;
        end else begin
          if (_T_16926) begin
            _T_16926 <= _T_16931;
          end
        end
      end else begin
        if (_T_16926) begin
          _T_16926 <= _T_16931;
        end
      end
    end
    if (reset) begin
      _T_16945_0 <= 1'h0;
    end else begin
      if (_T_17496) begin
        if (_T_17498) begin
          _T_16945_0 <= 1'h0;
        end else begin
          if (_T_17303) begin
            _T_16945_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_17303) begin
          _T_16945_0 <= 1'h1;
        end
      end
    end
    if (_T_17303) begin
      _T_16958_0 <= _T_530_0;
    end
    if (_T_542_0) begin
      if (5'h0 == _T_554_0) begin
        _T_17035_0_0 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h1 == _T_554_0) begin
        _T_17035_0_1 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h2 == _T_554_0) begin
        _T_17035_0_2 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h3 == _T_554_0) begin
        _T_17035_0_3 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h4 == _T_554_0) begin
        _T_17035_0_4 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h5 == _T_554_0) begin
        _T_17035_0_5 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h6 == _T_554_0) begin
        _T_17035_0_6 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h7 == _T_554_0) begin
        _T_17035_0_7 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h8 == _T_554_0) begin
        _T_17035_0_8 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h9 == _T_554_0) begin
        _T_17035_0_9 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'ha == _T_554_0) begin
        _T_17035_0_10 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'hb == _T_554_0) begin
        _T_17035_0_11 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'hc == _T_554_0) begin
        _T_17035_0_12 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'hd == _T_554_0) begin
        _T_17035_0_13 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'he == _T_554_0) begin
        _T_17035_0_14 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'hf == _T_554_0) begin
        _T_17035_0_15 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h10 == _T_554_0) begin
        _T_17035_0_16 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h11 == _T_554_0) begin
        _T_17035_0_17 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h12 == _T_554_0) begin
        _T_17035_0_18 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h13 == _T_554_0) begin
        _T_17035_0_19 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h14 == _T_554_0) begin
        _T_17035_0_20 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h15 == _T_554_0) begin
        _T_17035_0_21 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h16 == _T_554_0) begin
        _T_17035_0_22 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h17 == _T_554_0) begin
        _T_17035_0_23 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h18 == _T_554_0) begin
        _T_17035_0_24 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h19 == _T_554_0) begin
        _T_17035_0_25 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h1a == _T_554_0) begin
        _T_17035_0_26 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h1b == _T_554_0) begin
        _T_17035_0_27 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h1c == _T_554_0) begin
        _T_17035_0_28 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h1d == _T_554_0) begin
        _T_17035_0_29 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h1e == _T_554_0) begin
        _T_17035_0_30 <= _GEN_5;
      end
    end
    if (_T_542_0) begin
      if (5'h1f == _T_554_0) begin
        _T_17035_0_31 <= _GEN_5;
      end
    end
    if (reset) begin
      _T_17254_0 <= 1'h0;
    end else begin
      if (_T_17496) begin
        if (_T_17498) begin
          _T_17254_0 <= 1'h0;
        end else begin
          if (_T_17288) begin
            _T_17254_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_17288) begin
          _T_17254_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_17264 <= 1'h0;
    end else begin
      if (_T_17496) begin
        if (_T_17498) begin
          _T_17264 <= 1'h0;
        end else begin
          if (_T_17468) begin
            if (!(_T_17470)) begin
              _T_17264 <= _T_17474;
            end
          end
        end
      end else begin
        if (_T_17468) begin
          if (!(_T_17470)) begin
            _T_17264 <= _T_17474;
          end
        end
      end
    end
    if (reset) begin
      _T_17267 <= 1'h0;
    end else begin
      if (_T_17496) begin
        if (_T_17498) begin
          _T_17267 <= 1'h0;
        end else begin
          if (_T_17468) begin
            if (_T_17470) begin
              _T_17267 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_17468) begin
          if (_T_17470) begin
            _T_17267 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_17270 <= 1'h0;
    end else begin
      if (_T_17496) begin
        if (_T_17498) begin
          _T_17270 <= 1'h0;
        end else begin
          _T_17270 <= _T_17515;
        end
      end
    end
    if (reset) begin
      _T_17273 <= 1'h0;
    end else begin
      if (_T_17475) begin
        if (_T_17273) begin
          _T_17273 <= 1'h0;
        end else begin
          _T_17273 <= _T_17481;
        end
      end
    end
    if (reset) begin
      _T_17276 <= 1'h0;
    end else begin
      if (_T_17496) begin
        if (_T_17498) begin
          _T_17276 <= 1'h0;
        end else begin
          if (_T_17281) begin
            _T_17276 <= 1'h1;
          end
        end
      end else begin
        if (_T_17281) begin
          _T_17276 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_17534 <= 1'h0;
    end else begin
      if (_T_18104) begin
        if (_T_18106) begin
          _T_17534 <= 1'h0;
        end else begin
          if (_T_17534) begin
            _T_17534 <= _T_17539;
          end
        end
      end else begin
        if (_T_17534) begin
          _T_17534 <= _T_17539;
        end
      end
    end
    if (reset) begin
      _T_17553_0 <= 1'h0;
    end else begin
      if (_T_18104) begin
        if (_T_18106) begin
          _T_17553_0 <= 1'h0;
        end else begin
          if (_T_17911) begin
            _T_17553_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_17911) begin
          _T_17553_0 <= 1'h1;
        end
      end
    end
    if (_T_17911) begin
      _T_17566_0 <= _T_566_0;
    end
    if (_T_578_0) begin
      if (5'h0 == _T_590_0) begin
        _T_17643_0_0 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h1 == _T_590_0) begin
        _T_17643_0_1 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h2 == _T_590_0) begin
        _T_17643_0_2 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h3 == _T_590_0) begin
        _T_17643_0_3 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h4 == _T_590_0) begin
        _T_17643_0_4 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h5 == _T_590_0) begin
        _T_17643_0_5 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h6 == _T_590_0) begin
        _T_17643_0_6 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h7 == _T_590_0) begin
        _T_17643_0_7 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h8 == _T_590_0) begin
        _T_17643_0_8 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h9 == _T_590_0) begin
        _T_17643_0_9 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'ha == _T_590_0) begin
        _T_17643_0_10 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'hb == _T_590_0) begin
        _T_17643_0_11 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'hc == _T_590_0) begin
        _T_17643_0_12 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'hd == _T_590_0) begin
        _T_17643_0_13 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'he == _T_590_0) begin
        _T_17643_0_14 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'hf == _T_590_0) begin
        _T_17643_0_15 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h10 == _T_590_0) begin
        _T_17643_0_16 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h11 == _T_590_0) begin
        _T_17643_0_17 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h12 == _T_590_0) begin
        _T_17643_0_18 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h13 == _T_590_0) begin
        _T_17643_0_19 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h14 == _T_590_0) begin
        _T_17643_0_20 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h15 == _T_590_0) begin
        _T_17643_0_21 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h16 == _T_590_0) begin
        _T_17643_0_22 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h17 == _T_590_0) begin
        _T_17643_0_23 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h18 == _T_590_0) begin
        _T_17643_0_24 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h19 == _T_590_0) begin
        _T_17643_0_25 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h1a == _T_590_0) begin
        _T_17643_0_26 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h1b == _T_590_0) begin
        _T_17643_0_27 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h1c == _T_590_0) begin
        _T_17643_0_28 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h1d == _T_590_0) begin
        _T_17643_0_29 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h1e == _T_590_0) begin
        _T_17643_0_30 <= _GEN_6;
      end
    end
    if (_T_578_0) begin
      if (5'h1f == _T_590_0) begin
        _T_17643_0_31 <= _GEN_6;
      end
    end
    if (reset) begin
      _T_17862_0 <= 1'h0;
    end else begin
      if (_T_18104) begin
        if (_T_18106) begin
          _T_17862_0 <= 1'h0;
        end else begin
          if (_T_17896) begin
            _T_17862_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_17896) begin
          _T_17862_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_17872 <= 1'h0;
    end else begin
      if (_T_18104) begin
        if (_T_18106) begin
          _T_17872 <= 1'h0;
        end else begin
          if (_T_18076) begin
            if (!(_T_18078)) begin
              _T_17872 <= _T_18082;
            end
          end
        end
      end else begin
        if (_T_18076) begin
          if (!(_T_18078)) begin
            _T_17872 <= _T_18082;
          end
        end
      end
    end
    if (reset) begin
      _T_17875 <= 1'h0;
    end else begin
      if (_T_18104) begin
        if (_T_18106) begin
          _T_17875 <= 1'h0;
        end else begin
          if (_T_18076) begin
            if (_T_18078) begin
              _T_17875 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_18076) begin
          if (_T_18078) begin
            _T_17875 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_17878 <= 1'h0;
    end else begin
      if (_T_18104) begin
        if (_T_18106) begin
          _T_17878 <= 1'h0;
        end else begin
          _T_17878 <= _T_18123;
        end
      end
    end
    if (reset) begin
      _T_17881 <= 1'h0;
    end else begin
      if (_T_18083) begin
        if (_T_17881) begin
          _T_17881 <= 1'h0;
        end else begin
          _T_17881 <= _T_18089;
        end
      end
    end
    if (reset) begin
      _T_17884 <= 1'h0;
    end else begin
      if (_T_18104) begin
        if (_T_18106) begin
          _T_17884 <= 1'h0;
        end else begin
          if (_T_17889) begin
            _T_17884 <= 1'h1;
          end
        end
      end else begin
        if (_T_17889) begin
          _T_17884 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_18142 <= 1'h0;
    end else begin
      if (_T_18712) begin
        if (_T_18714) begin
          _T_18142 <= 1'h0;
        end else begin
          if (_T_18142) begin
            _T_18142 <= _T_18147;
          end
        end
      end else begin
        if (_T_18142) begin
          _T_18142 <= _T_18147;
        end
      end
    end
    if (reset) begin
      _T_18161_0 <= 1'h0;
    end else begin
      if (_T_18712) begin
        if (_T_18714) begin
          _T_18161_0 <= 1'h0;
        end else begin
          if (_T_18519) begin
            _T_18161_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_18519) begin
          _T_18161_0 <= 1'h1;
        end
      end
    end
    if (_T_18519) begin
      _T_18174_0 <= _T_602_0;
    end
    if (_T_614_0) begin
      if (5'h0 == _T_626_0) begin
        _T_18251_0_0 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h1 == _T_626_0) begin
        _T_18251_0_1 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h2 == _T_626_0) begin
        _T_18251_0_2 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h3 == _T_626_0) begin
        _T_18251_0_3 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h4 == _T_626_0) begin
        _T_18251_0_4 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h5 == _T_626_0) begin
        _T_18251_0_5 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h6 == _T_626_0) begin
        _T_18251_0_6 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h7 == _T_626_0) begin
        _T_18251_0_7 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h8 == _T_626_0) begin
        _T_18251_0_8 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h9 == _T_626_0) begin
        _T_18251_0_9 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'ha == _T_626_0) begin
        _T_18251_0_10 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'hb == _T_626_0) begin
        _T_18251_0_11 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'hc == _T_626_0) begin
        _T_18251_0_12 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'hd == _T_626_0) begin
        _T_18251_0_13 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'he == _T_626_0) begin
        _T_18251_0_14 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'hf == _T_626_0) begin
        _T_18251_0_15 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h10 == _T_626_0) begin
        _T_18251_0_16 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h11 == _T_626_0) begin
        _T_18251_0_17 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h12 == _T_626_0) begin
        _T_18251_0_18 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h13 == _T_626_0) begin
        _T_18251_0_19 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h14 == _T_626_0) begin
        _T_18251_0_20 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h15 == _T_626_0) begin
        _T_18251_0_21 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h16 == _T_626_0) begin
        _T_18251_0_22 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h17 == _T_626_0) begin
        _T_18251_0_23 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h18 == _T_626_0) begin
        _T_18251_0_24 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h19 == _T_626_0) begin
        _T_18251_0_25 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h1a == _T_626_0) begin
        _T_18251_0_26 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h1b == _T_626_0) begin
        _T_18251_0_27 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h1c == _T_626_0) begin
        _T_18251_0_28 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h1d == _T_626_0) begin
        _T_18251_0_29 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h1e == _T_626_0) begin
        _T_18251_0_30 <= _GEN_7;
      end
    end
    if (_T_614_0) begin
      if (5'h1f == _T_626_0) begin
        _T_18251_0_31 <= _GEN_7;
      end
    end
    if (reset) begin
      _T_18470_0 <= 1'h0;
    end else begin
      if (_T_18712) begin
        if (_T_18714) begin
          _T_18470_0 <= 1'h0;
        end else begin
          if (_T_18504) begin
            _T_18470_0 <= 1'h1;
          end
        end
      end else begin
        if (_T_18504) begin
          _T_18470_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_18480 <= 1'h0;
    end else begin
      if (_T_18712) begin
        if (_T_18714) begin
          _T_18480 <= 1'h0;
        end else begin
          if (_T_18684) begin
            if (!(_T_18686)) begin
              _T_18480 <= _T_18690;
            end
          end
        end
      end else begin
        if (_T_18684) begin
          if (!(_T_18686)) begin
            _T_18480 <= _T_18690;
          end
        end
      end
    end
    if (reset) begin
      _T_18483 <= 1'h0;
    end else begin
      if (_T_18712) begin
        if (_T_18714) begin
          _T_18483 <= 1'h0;
        end else begin
          if (_T_18684) begin
            if (_T_18686) begin
              _T_18483 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_18684) begin
          if (_T_18686) begin
            _T_18483 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_18486 <= 1'h0;
    end else begin
      if (_T_18712) begin
        if (_T_18714) begin
          _T_18486 <= 1'h0;
        end else begin
          _T_18486 <= _T_18731;
        end
      end
    end
    if (reset) begin
      _T_18489 <= 1'h0;
    end else begin
      if (_T_18691) begin
        if (_T_18489) begin
          _T_18489 <= 1'h0;
        end else begin
          _T_18489 <= _T_18697;
        end
      end
    end
    if (reset) begin
      _T_18492 <= 1'h0;
    end else begin
      if (_T_18712) begin
        if (_T_18714) begin
          _T_18492 <= 1'h0;
        end else begin
          if (_T_18497) begin
            _T_18492 <= 1'h1;
          end
        end
      end else begin
        if (_T_18497) begin
          _T_18492 <= 1'h1;
        end
      end
    end
  end
endmodule
module PassThrough(
  input        clock,
  input        reset,
  input  [7:0] io_inputWord,
  input        io_inputValid,
  input        io_inputFinished,
  output       io_inputReady,
  output [7:0] io_outputWord,
  output       io_outputValid,
  output       io_outputFinished,
  input        io_outputReady
);
  reg [7:0] _T_11;
  reg [31:0] _RAND_0;
  reg  _T_14;
  reg [31:0] _RAND_1;
  reg  _T_17;
  reg [31:0] _RAND_2;
  wire  _T_21;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  reg  _T_31;
  reg [31:0] _RAND_3;
  wire  _T_35;
  wire  _T_37;
  wire  _T_38;
  wire  _T_41;
  wire  _T_45;
  wire  _T_46;
  wire [1:0] _T_48;
  wire  _T_49;
  wire  _GEN_0;
  wire  _T_55;
  wire  _T_56;
  wire  _T_57;
  wire [7:0] _GEN_1;
  wire  _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire  _T_67;
  wire [7:0] _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire [7:0] _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _T_86;
  wire  _T_91;
  assign _T_23 = io_outputValid == 1'h0;
  assign _T_24 = _T_23 | io_outputReady;
  assign _T_25 = _T_21 & _T_24;
  assign _T_35 = _T_31 == 1'h0;
  assign _T_37 = _T_14 == 1'h0;
  assign _T_38 = _T_35 & _T_37;
  assign _T_41 = _T_38 | _T_25;
  assign _T_45 = _T_21 == 1'h0;
  assign _T_46 = _T_31 & _T_45;
  assign _T_48 = _T_31 + 1'h1;
  assign _T_49 = _T_48[0:0];
  assign _GEN_0 = _T_46 ? _T_49 : _T_31;
  assign _T_55 = _T_17 == 1'h0;
  assign _T_56 = io_inputFinished & _T_55;
  assign _T_57 = _T_56 | io_inputValid;
  assign _GEN_1 = _T_37 ? io_inputWord : _T_11;
  assign _GEN_2 = _T_37 ? io_inputFinished : _T_17;
  assign _GEN_3 = _T_37 ? _T_57 : _T_14;
  assign _GEN_4 = _T_37 ? _T_57 : 1'h1;
  assign _GEN_10 = _T_25 ? io_inputWord : _T_11;
  assign _GEN_11 = _T_25 ? io_inputFinished : _T_17;
  assign _GEN_12 = _T_25 ? _T_57 : _T_14;
  assign _GEN_13 = _T_25 ? _T_67 : _GEN_0;
  assign _GEN_14 = _T_35 ? _GEN_1 : _GEN_10;
  assign _GEN_15 = _T_35 ? _GEN_2 : _GEN_11;
  assign _GEN_16 = _T_35 ? _GEN_3 : _GEN_12;
  assign _GEN_17 = _T_35 ? _GEN_4 : _GEN_13;
  assign _T_86 = _T_17 & _T_35;
  assign _T_91 = _T_21 & _T_55;
  assign io_inputReady = _T_41;
  assign io_outputWord = _T_11;
  assign io_outputValid = _T_91;
  assign io_outputFinished = _T_86;
  assign _T_21 = _T_31;
  assign _T_67 = _T_57;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_11 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_14 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_17 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_31 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_35) begin
      if (_T_37) begin
        _T_11 <= io_inputWord;
      end
    end else begin
      if (_T_25) begin
        _T_11 <= io_inputWord;
      end
    end
    if (reset) begin
      _T_14 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_37) begin
          _T_14 <= _T_57;
        end
      end else begin
        if (_T_25) begin
          _T_14 <= _T_57;
        end
      end
    end
    if (reset) begin
      _T_17 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_37) begin
          _T_17 <= io_inputFinished;
        end
      end else begin
        if (_T_25) begin
          _T_17 <= io_inputFinished;
        end
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_37) begin
          _T_31 <= _T_57;
        end else begin
          _T_31 <= 1'h1;
        end
      end else begin
        if (_T_25) begin
          _T_31 <= _T_67;
        end else begin
          if (_T_46) begin
            _T_31 <= _T_49;
          end
        end
      end
    end
  end
endmodule
module DualPortBRAM(
  input         clock,
  input  [4:0]  io_a_addr,
  input  [31:0] io_a_din,
  input         io_a_wr,
  input  [4:0]  io_b_addr,
  output [31:0] io_b_dout
);
  reg [31:0] mem [0:31];
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_16_data;
  wire [4:0] mem__T_16_addr;
  wire [31:0] mem__T_22_data;
  wire [4:0] mem__T_22_addr;
  wire [31:0] mem__T_17_data;
  wire [4:0] mem__T_17_addr;
  wire  mem__T_17_mask;
  wire  mem__T_17_en;
  wire [31:0] mem__T_23_data;
  wire [4:0] mem__T_23_addr;
  wire  mem__T_23_mask;
  wire  mem__T_23_en;
  reg [4:0] regAddrA;
  reg [31:0] _RAND_1;
  reg [4:0] regAddrB;
  reg [31:0] _RAND_2;
  assign mem__T_16_addr = regAddrA;
  assign mem__T_16_data = mem[mem__T_16_addr];
  assign mem__T_22_addr = regAddrB;
  assign mem__T_22_data = mem[mem__T_22_addr];
  assign mem__T_17_data = io_a_din;
  assign mem__T_17_addr = io_a_addr;
  assign mem__T_17_mask = io_a_wr;
  assign mem__T_17_en = io_a_wr;
  assign mem__T_23_data = 32'h0;
  assign mem__T_23_addr = io_b_addr;
  assign mem__T_23_mask = 1'h0;
  assign mem__T_23_en = 1'h0;
  assign io_b_dout = mem__T_22_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  regAddrA = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  regAddrB = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_17_en & mem__T_17_mask) begin
      mem[mem__T_17_addr] <= mem__T_17_data;
    end
    if(mem__T_23_en & mem__T_23_mask) begin
      mem[mem__T_23_addr] <= mem__T_23_data;
    end
    regAddrA <= io_a_addr;
    regAddrB <= io_b_addr;
  end
endmodule
module InnerCore(
  input         clock,
  input         reset,
  input  [31:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  input  [10:0] io_inputBits,
  output        io_inputMemConsumed,
  input         io_inputFinished,
  output [31:0] io_outputMemBlock,
  output        io_outputMemBlockValid,
  input         io_outputMemBlockReady,
  output [10:0] io_outputBits,
  output        io_outputFinished
);
  wire  inner_clock;
  wire  inner_reset;
  wire [7:0] inner_io_inputWord;
  wire  inner_io_inputValid;
  wire  inner_io_inputFinished;
  wire  inner_io_inputReady;
  wire [7:0] inner_io_outputWord;
  wire  inner_io_outputValid;
  wire  inner_io_outputFinished;
  wire  inner_io_outputReady;
  reg  inputMemBlock_0;
  reg [31:0] _RAND_0;
  reg  inputMemBlock_1;
  reg [31:0] _RAND_1;
  reg  inputMemBlock_2;
  reg [31:0] _RAND_2;
  reg  inputMemBlock_3;
  reg [31:0] _RAND_3;
  reg  inputMemBlock_4;
  reg [31:0] _RAND_4;
  reg  inputMemBlock_5;
  reg [31:0] _RAND_5;
  reg  inputMemBlock_6;
  reg [31:0] _RAND_6;
  reg  inputMemBlock_7;
  reg [31:0] _RAND_7;
  reg  inputMemBlock_8;
  reg [31:0] _RAND_8;
  reg  inputMemBlock_9;
  reg [31:0] _RAND_9;
  reg  inputMemBlock_10;
  reg [31:0] _RAND_10;
  reg  inputMemBlock_11;
  reg [31:0] _RAND_11;
  reg  inputMemBlock_12;
  reg [31:0] _RAND_12;
  reg  inputMemBlock_13;
  reg [31:0] _RAND_13;
  reg  inputMemBlock_14;
  reg [31:0] _RAND_14;
  reg  inputMemBlock_15;
  reg [31:0] _RAND_15;
  reg  inputMemBlock_16;
  reg [31:0] _RAND_16;
  reg  inputMemBlock_17;
  reg [31:0] _RAND_17;
  reg  inputMemBlock_18;
  reg [31:0] _RAND_18;
  reg  inputMemBlock_19;
  reg [31:0] _RAND_19;
  reg  inputMemBlock_20;
  reg [31:0] _RAND_20;
  reg  inputMemBlock_21;
  reg [31:0] _RAND_21;
  reg  inputMemBlock_22;
  reg [31:0] _RAND_22;
  reg  inputMemBlock_23;
  reg [31:0] _RAND_23;
  reg  inputMemBlock_24;
  reg [31:0] _RAND_24;
  reg  inputMemBlock_25;
  reg [31:0] _RAND_25;
  reg  inputMemBlock_26;
  reg [31:0] _RAND_26;
  reg  inputMemBlock_27;
  reg [31:0] _RAND_27;
  reg  inputMemBlock_28;
  reg [31:0] _RAND_28;
  reg  inputMemBlock_29;
  reg [31:0] _RAND_29;
  reg  inputMemBlock_30;
  reg [31:0] _RAND_30;
  reg  inputMemBlock_31;
  reg [31:0] _RAND_31;
  reg [5:0] inputPieceBitsRemaining;
  reg [31:0] _RAND_32;
  reg [10:0] inputBitsRemaining;
  reg [31:0] _RAND_33;
  reg  outputMemBlock_0;
  reg [31:0] _RAND_34;
  reg  outputMemBlock_1;
  reg [31:0] _RAND_35;
  reg  outputMemBlock_2;
  reg [31:0] _RAND_36;
  reg  outputMemBlock_3;
  reg [31:0] _RAND_37;
  reg  outputMemBlock_4;
  reg [31:0] _RAND_38;
  reg  outputMemBlock_5;
  reg [31:0] _RAND_39;
  reg  outputMemBlock_6;
  reg [31:0] _RAND_40;
  reg  outputMemBlock_7;
  reg [31:0] _RAND_41;
  reg  outputMemBlock_8;
  reg [31:0] _RAND_42;
  reg  outputMemBlock_9;
  reg [31:0] _RAND_43;
  reg  outputMemBlock_10;
  reg [31:0] _RAND_44;
  reg  outputMemBlock_11;
  reg [31:0] _RAND_45;
  reg  outputMemBlock_12;
  reg [31:0] _RAND_46;
  reg  outputMemBlock_13;
  reg [31:0] _RAND_47;
  reg  outputMemBlock_14;
  reg [31:0] _RAND_48;
  reg  outputMemBlock_15;
  reg [31:0] _RAND_49;
  reg  outputMemBlock_16;
  reg [31:0] _RAND_50;
  reg  outputMemBlock_17;
  reg [31:0] _RAND_51;
  reg  outputMemBlock_18;
  reg [31:0] _RAND_52;
  reg  outputMemBlock_19;
  reg [31:0] _RAND_53;
  reg  outputMemBlock_20;
  reg [31:0] _RAND_54;
  reg  outputMemBlock_21;
  reg [31:0] _RAND_55;
  reg  outputMemBlock_22;
  reg [31:0] _RAND_56;
  reg  outputMemBlock_23;
  reg [31:0] _RAND_57;
  reg  outputMemBlock_24;
  reg [31:0] _RAND_58;
  reg  outputMemBlock_25;
  reg [31:0] _RAND_59;
  reg  outputMemBlock_26;
  reg [31:0] _RAND_60;
  reg  outputMemBlock_27;
  reg [31:0] _RAND_61;
  reg  outputMemBlock_28;
  reg [31:0] _RAND_62;
  reg  outputMemBlock_29;
  reg [31:0] _RAND_63;
  reg  outputMemBlock_30;
  reg [31:0] _RAND_64;
  reg  outputMemBlock_31;
  reg [31:0] _RAND_65;
  reg [10:0] outputBits;
  reg [31:0] _RAND_66;
  reg [5:0] outputPieceBits;
  reg [31:0] _RAND_67;
  wire  inputBram_clock;
  wire [4:0] inputBram_io_a_addr;
  wire [31:0] inputBram_io_a_din;
  wire  inputBram_io_a_wr;
  wire [4:0] inputBram_io_b_addr;
  wire [31:0] inputBram_io_b_dout;
  reg [4:0] inputReadAddr;
  reg [31:0] _RAND_68;
  wire  outputBram_clock;
  wire [4:0] outputBram_io_a_addr;
  wire [31:0] outputBram_io_a_din;
  wire  outputBram_io_a_wr;
  wire [4:0] outputBram_io_b_addr;
  wire [31:0] outputBram_io_b_dout;
  reg [4:0] outputWriteAddr;
  reg [31:0] _RAND_69;
  reg [4:0] outputReadAddr;
  reg [31:0] _RAND_70;
  wire  _T_102;
  wire  _T_103;
  wire [10:0] _GEN_0;
  wire [4:0] inputReadAddrFinal;
  wire  _T_107;
  wire  _T_109;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire [6:0] _T_115;
  wire [6:0] _T_116;
  wire [5:0] _T_117;
  wire  _T_119;
  wire  _T_120;
  wire  _T_121;
  wire [11:0] _T_125;
  wire [11:0] _T_126;
  wire [10:0] _T_127;
  wire [10:0] _T_128;
  wire  _T_130;
  wire [10:0] _T_132;
  wire  _T_134;
  wire [5:0] _T_136;
  wire [4:0] _T_137;
  wire [4:0] _T_138;
  wire  _T_142;
  wire  _T_143;
  wire  _T_144;
  wire  _T_145;
  wire  _T_146;
  wire  _T_147;
  wire  _T_148;
  wire  _T_149;
  wire  _T_150;
  wire  _T_151;
  wire  _T_152;
  wire  _T_153;
  wire  _T_154;
  wire  _T_155;
  wire  _T_156;
  wire  _T_157;
  wire  _T_158;
  wire  _T_159;
  wire  _T_160;
  wire  _T_161;
  wire  _T_162;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _T_166;
  wire  _T_167;
  wire  _T_168;
  wire  _T_169;
  wire  _T_170;
  wire  _T_171;
  wire  _T_172;
  wire  _T_173;
  wire [10:0] _GEN_1;
  wire [10:0] _GEN_2;
  wire [4:0] _GEN_3;
  wire [4:0] _GEN_4;
  wire  _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _T_182;
  wire  _T_183;
  wire [10:0] _GEN_37;
  wire [10:0] _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire  _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire [1:0] _T_192;
  wire [1:0] _T_193;
  wire [3:0] _T_194;
  wire [1:0] _T_195;
  wire [1:0] _T_196;
  wire [3:0] _T_197;
  wire [7:0] _T_198;
  wire [1:0] _T_199;
  wire [1:0] _T_200;
  wire [3:0] _T_201;
  wire [1:0] _T_202;
  wire [1:0] _T_203;
  wire [3:0] _T_204;
  wire [7:0] _T_205;
  wire [15:0] _T_206;
  wire [1:0] _T_207;
  wire [1:0] _T_208;
  wire [3:0] _T_209;
  wire [1:0] _T_210;
  wire [1:0] _T_211;
  wire [3:0] _T_212;
  wire [7:0] _T_213;
  wire [1:0] _T_214;
  wire [1:0] _T_215;
  wire [3:0] _T_216;
  wire [1:0] _T_217;
  wire [1:0] _T_218;
  wire [3:0] _T_219;
  wire [7:0] _T_220;
  wire [15:0] _T_221;
  wire [31:0] _T_222;
  wire [7:0] nextWord;
  wire  _T_226;
  wire  _T_229;
  wire  _T_231;
  wire  _T_233;
  wire  _T_234;
  wire  _T_236;
  wire  _T_237;
  wire  _T_239;
  wire  _T_240;
  wire  _T_241;
  wire  _T_242;
  wire  _T_243;
  wire  _T_244;
  wire  _T_245;
  wire  _T_246;
  wire  _T_247;
  wire  _T_248;
  wire  _T_249;
  wire  _T_251;
  wire [6:0] _T_254;
  wire [5:0] _T_255;
  wire [5:0] _T_256;
  wire [5:0] _T_260;
  wire [4:0] _T_261;
  wire [4:0] _T_262;
  wire [11:0] _T_264;
  wire [10:0] _T_265;
  wire [10:0] _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_76;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire  _GEN_83;
  wire  _GEN_84;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire  _GEN_90;
  wire  _GEN_91;
  wire  _GEN_92;
  wire  _GEN_93;
  wire  _GEN_94;
  wire  _GEN_95;
  wire [5:0] _GEN_96;
  wire [4:0] _GEN_97;
  wire [10:0] _GEN_98;
  wire [1:0] _T_268;
  wire [1:0] _T_269;
  wire [3:0] _T_270;
  wire [1:0] _T_271;
  wire [1:0] _T_272;
  wire [3:0] _T_273;
  wire [7:0] _T_274;
  wire [1:0] _T_275;
  wire [1:0] _T_276;
  wire [3:0] _T_277;
  wire [1:0] _T_278;
  wire [1:0] _T_279;
  wire [3:0] _T_280;
  wire [7:0] _T_281;
  wire [15:0] _T_282;
  wire [1:0] _T_283;
  wire [1:0] _T_284;
  wire [3:0] _T_285;
  wire [1:0] _T_286;
  wire [1:0] _T_287;
  wire [3:0] _T_288;
  wire [7:0] _T_289;
  wire [1:0] _T_290;
  wire [1:0] _T_291;
  wire [3:0] _T_292;
  wire [1:0] _T_293;
  wire [1:0] _T_294;
  wire [3:0] _T_295;
  wire [7:0] _T_296;
  wire [15:0] _T_297;
  wire [31:0] _T_298;
  reg  outputReadingStartedPrev;
  reg [31:0] _RAND_71;
  reg  outputReadingStarted;
  reg [31:0] _RAND_72;
  wire  _T_305;
  wire  _T_309;
  wire  _T_310;
  wire  _T_313;
  wire  _T_314;
  wire  _T_315;
  wire  _GEN_99;
  wire  _T_318;
  wire  _T_319;
  wire  _GEN_100;
  wire  _T_321;
  wire  _T_323;
  wire  _T_325;
  wire  _T_326;
  wire [5:0] _T_328;
  wire [4:0] _T_329;
  wire  _T_331;
  wire [10:0] _GEN_101;
  wire [4:0] _GEN_102;
  wire [10:0] _GEN_103;
  wire  _T_336;
  wire  _T_337;
  wire  _T_340;
  wire  _T_343;
  wire  _GEN_104;
  wire  _GEN_105;
  wire [4:0] _GEN_106;
  PassThrough inner (
    .clock(inner_clock),
    .reset(inner_reset),
    .io_inputWord(inner_io_inputWord),
    .io_inputValid(inner_io_inputValid),
    .io_inputFinished(inner_io_inputFinished),
    .io_inputReady(inner_io_inputReady),
    .io_outputWord(inner_io_outputWord),
    .io_outputValid(inner_io_outputValid),
    .io_outputFinished(inner_io_outputFinished),
    .io_outputReady(inner_io_outputReady)
  );
  DualPortBRAM inputBram (
    .clock(inputBram_clock),
    .io_a_addr(inputBram_io_a_addr),
    .io_a_din(inputBram_io_a_din),
    .io_a_wr(inputBram_io_a_wr),
    .io_b_addr(inputBram_io_b_addr),
    .io_b_dout(inputBram_io_b_dout)
  );
  DualPortBRAM outputBram (
    .clock(outputBram_clock),
    .io_a_addr(outputBram_io_a_addr),
    .io_a_din(outputBram_io_a_din),
    .io_a_wr(outputBram_io_a_wr),
    .io_b_addr(outputBram_io_b_addr),
    .io_b_dout(outputBram_io_b_dout)
  );
  assign _T_102 = io_inputMemIdx == 5'h1;
  assign _T_103 = io_inputMemBlockValid & _T_102;
  assign _GEN_0 = _T_103 ? io_inputBits : inputBitsRemaining;
  assign _T_107 = inputPieceBitsRemaining == 6'h0;
  assign _T_109 = inputBitsRemaining == 11'h0;
  assign _T_111 = _T_109 == 1'h0;
  assign _T_112 = _T_107 & _T_111;
  assign _T_113 = inner_io_inputValid & inner_io_inputReady;
  assign _T_115 = inputPieceBitsRemaining - 6'h8;
  assign _T_116 = $unsigned(_T_115);
  assign _T_117 = _T_116[5:0];
  assign _T_119 = _T_117 == 6'h0;
  assign _T_120 = _T_113 & _T_119;
  assign _T_121 = _T_112 | _T_120;
  assign _T_125 = inputBitsRemaining - 11'h8;
  assign _T_126 = $unsigned(_T_125);
  assign _T_127 = _T_126[10:0];
  assign _T_128 = _T_107 ? inputBitsRemaining : _T_127;
  assign _T_130 = _T_128 < 11'h20;
  assign _T_132 = _T_130 ? _T_128 : 11'h20;
  assign _T_134 = _T_128 == 11'h0;
  assign _T_136 = inputReadAddr + 5'h1;
  assign _T_137 = _T_136[4:0];
  assign _T_138 = _T_134 ? inputReadAddr : _T_137;
  assign _T_142 = inputBram_io_b_dout[0];
  assign _T_143 = inputBram_io_b_dout[1];
  assign _T_144 = inputBram_io_b_dout[2];
  assign _T_145 = inputBram_io_b_dout[3];
  assign _T_146 = inputBram_io_b_dout[4];
  assign _T_147 = inputBram_io_b_dout[5];
  assign _T_148 = inputBram_io_b_dout[6];
  assign _T_149 = inputBram_io_b_dout[7];
  assign _T_150 = inputBram_io_b_dout[8];
  assign _T_151 = inputBram_io_b_dout[9];
  assign _T_152 = inputBram_io_b_dout[10];
  assign _T_153 = inputBram_io_b_dout[11];
  assign _T_154 = inputBram_io_b_dout[12];
  assign _T_155 = inputBram_io_b_dout[13];
  assign _T_156 = inputBram_io_b_dout[14];
  assign _T_157 = inputBram_io_b_dout[15];
  assign _T_158 = inputBram_io_b_dout[16];
  assign _T_159 = inputBram_io_b_dout[17];
  assign _T_160 = inputBram_io_b_dout[18];
  assign _T_161 = inputBram_io_b_dout[19];
  assign _T_162 = inputBram_io_b_dout[20];
  assign _T_163 = inputBram_io_b_dout[21];
  assign _T_164 = inputBram_io_b_dout[22];
  assign _T_165 = inputBram_io_b_dout[23];
  assign _T_166 = inputBram_io_b_dout[24];
  assign _T_167 = inputBram_io_b_dout[25];
  assign _T_168 = inputBram_io_b_dout[26];
  assign _T_169 = inputBram_io_b_dout[27];
  assign _T_170 = inputBram_io_b_dout[28];
  assign _T_171 = inputBram_io_b_dout[29];
  assign _T_172 = inputBram_io_b_dout[30];
  assign _T_173 = inputBram_io_b_dout[31];
  assign _GEN_1 = _T_121 ? _T_132 : {{5'd0}, inputPieceBitsRemaining};
  assign _GEN_2 = _T_121 ? _T_128 : _GEN_0;
  assign _GEN_3 = _T_121 ? _T_138 : inputReadAddr;
  assign _GEN_4 = _T_121 ? _T_137 : inputReadAddr;
  assign _GEN_5 = _T_121 ? _T_142 : inputMemBlock_0;
  assign _GEN_6 = _T_121 ? _T_143 : inputMemBlock_1;
  assign _GEN_7 = _T_121 ? _T_144 : inputMemBlock_2;
  assign _GEN_8 = _T_121 ? _T_145 : inputMemBlock_3;
  assign _GEN_9 = _T_121 ? _T_146 : inputMemBlock_4;
  assign _GEN_10 = _T_121 ? _T_147 : inputMemBlock_5;
  assign _GEN_11 = _T_121 ? _T_148 : inputMemBlock_6;
  assign _GEN_12 = _T_121 ? _T_149 : inputMemBlock_7;
  assign _GEN_13 = _T_121 ? _T_150 : inputMemBlock_8;
  assign _GEN_14 = _T_121 ? _T_151 : inputMemBlock_9;
  assign _GEN_15 = _T_121 ? _T_152 : inputMemBlock_10;
  assign _GEN_16 = _T_121 ? _T_153 : inputMemBlock_11;
  assign _GEN_17 = _T_121 ? _T_154 : inputMemBlock_12;
  assign _GEN_18 = _T_121 ? _T_155 : inputMemBlock_13;
  assign _GEN_19 = _T_121 ? _T_156 : inputMemBlock_14;
  assign _GEN_20 = _T_121 ? _T_157 : inputMemBlock_15;
  assign _GEN_21 = _T_121 ? _T_158 : inputMemBlock_16;
  assign _GEN_22 = _T_121 ? _T_159 : inputMemBlock_17;
  assign _GEN_23 = _T_121 ? _T_160 : inputMemBlock_18;
  assign _GEN_24 = _T_121 ? _T_161 : inputMemBlock_19;
  assign _GEN_25 = _T_121 ? _T_162 : inputMemBlock_20;
  assign _GEN_26 = _T_121 ? _T_163 : inputMemBlock_21;
  assign _GEN_27 = _T_121 ? _T_164 : inputMemBlock_22;
  assign _GEN_28 = _T_121 ? _T_165 : inputMemBlock_23;
  assign _GEN_29 = _T_121 ? _T_166 : inputMemBlock_24;
  assign _GEN_30 = _T_121 ? _T_167 : inputMemBlock_25;
  assign _GEN_31 = _T_121 ? _T_168 : inputMemBlock_26;
  assign _GEN_32 = _T_121 ? _T_169 : inputMemBlock_27;
  assign _GEN_33 = _T_121 ? _T_170 : inputMemBlock_28;
  assign _GEN_34 = _T_121 ? _T_171 : inputMemBlock_29;
  assign _GEN_35 = _T_121 ? _T_172 : inputMemBlock_30;
  assign _GEN_36 = _T_121 ? _T_173 : inputMemBlock_31;
  assign _T_182 = _T_119 == 1'h0;
  assign _T_183 = _T_113 & _T_182;
  assign _GEN_37 = _T_183 ? {{5'd0}, _T_117} : _GEN_1;
  assign _GEN_38 = _T_183 ? _T_127 : _GEN_2;
  assign _GEN_39 = _T_183 ? inputMemBlock_8 : _GEN_5;
  assign _GEN_40 = _T_183 ? inputMemBlock_9 : _GEN_6;
  assign _GEN_41 = _T_183 ? inputMemBlock_10 : _GEN_7;
  assign _GEN_42 = _T_183 ? inputMemBlock_11 : _GEN_8;
  assign _GEN_43 = _T_183 ? inputMemBlock_12 : _GEN_9;
  assign _GEN_44 = _T_183 ? inputMemBlock_13 : _GEN_10;
  assign _GEN_45 = _T_183 ? inputMemBlock_14 : _GEN_11;
  assign _GEN_46 = _T_183 ? inputMemBlock_15 : _GEN_12;
  assign _GEN_47 = _T_183 ? inputMemBlock_16 : _GEN_13;
  assign _GEN_48 = _T_183 ? inputMemBlock_17 : _GEN_14;
  assign _GEN_49 = _T_183 ? inputMemBlock_18 : _GEN_15;
  assign _GEN_50 = _T_183 ? inputMemBlock_19 : _GEN_16;
  assign _GEN_51 = _T_183 ? inputMemBlock_20 : _GEN_17;
  assign _GEN_52 = _T_183 ? inputMemBlock_21 : _GEN_18;
  assign _GEN_53 = _T_183 ? inputMemBlock_22 : _GEN_19;
  assign _GEN_54 = _T_183 ? inputMemBlock_23 : _GEN_20;
  assign _GEN_55 = _T_183 ? inputMemBlock_24 : _GEN_21;
  assign _GEN_56 = _T_183 ? inputMemBlock_25 : _GEN_22;
  assign _GEN_57 = _T_183 ? inputMemBlock_26 : _GEN_23;
  assign _GEN_58 = _T_183 ? inputMemBlock_27 : _GEN_24;
  assign _GEN_59 = _T_183 ? inputMemBlock_28 : _GEN_25;
  assign _GEN_60 = _T_183 ? inputMemBlock_29 : _GEN_26;
  assign _GEN_61 = _T_183 ? inputMemBlock_30 : _GEN_27;
  assign _GEN_62 = _T_183 ? inputMemBlock_31 : _GEN_28;
  assign _T_192 = {inputMemBlock_1,inputMemBlock_0};
  assign _T_193 = {inputMemBlock_3,inputMemBlock_2};
  assign _T_194 = {_T_193,_T_192};
  assign _T_195 = {inputMemBlock_5,inputMemBlock_4};
  assign _T_196 = {inputMemBlock_7,inputMemBlock_6};
  assign _T_197 = {_T_196,_T_195};
  assign _T_198 = {_T_197,_T_194};
  assign _T_199 = {inputMemBlock_9,inputMemBlock_8};
  assign _T_200 = {inputMemBlock_11,inputMemBlock_10};
  assign _T_201 = {_T_200,_T_199};
  assign _T_202 = {inputMemBlock_13,inputMemBlock_12};
  assign _T_203 = {inputMemBlock_15,inputMemBlock_14};
  assign _T_204 = {_T_203,_T_202};
  assign _T_205 = {_T_204,_T_201};
  assign _T_206 = {_T_205,_T_198};
  assign _T_207 = {inputMemBlock_17,inputMemBlock_16};
  assign _T_208 = {inputMemBlock_19,inputMemBlock_18};
  assign _T_209 = {_T_208,_T_207};
  assign _T_210 = {inputMemBlock_21,inputMemBlock_20};
  assign _T_211 = {inputMemBlock_23,inputMemBlock_22};
  assign _T_212 = {_T_211,_T_210};
  assign _T_213 = {_T_212,_T_209};
  assign _T_214 = {inputMemBlock_25,inputMemBlock_24};
  assign _T_215 = {inputMemBlock_27,inputMemBlock_26};
  assign _T_216 = {_T_215,_T_214};
  assign _T_217 = {inputMemBlock_29,inputMemBlock_28};
  assign _T_218 = {inputMemBlock_31,inputMemBlock_30};
  assign _T_219 = {_T_218,_T_217};
  assign _T_220 = {_T_219,_T_216};
  assign _T_221 = {_T_220,_T_213};
  assign _T_222 = {_T_221,_T_206};
  assign nextWord = _T_222[7:0];
  assign _T_226 = _T_107 == 1'h0;
  assign _T_229 = io_inputFinished & _T_109;
  assign _T_231 = outputBits == 11'h400;
  assign _T_233 = _T_231 == 1'h0;
  assign _T_234 = inner_io_outputValid & inner_io_outputReady;
  assign _T_236 = outputPieceBits > 6'h0;
  assign _T_237 = inner_io_outputFinished & _T_236;
  assign _T_239 = outputPieceBits < 6'h20;
  assign _T_240 = _T_237 & _T_239;
  assign _T_241 = _T_234 | _T_240;
  assign _T_242 = inner_io_outputWord[7];
  assign _T_243 = inner_io_outputWord[6];
  assign _T_244 = inner_io_outputWord[5];
  assign _T_245 = inner_io_outputWord[4];
  assign _T_246 = inner_io_outputWord[3];
  assign _T_247 = inner_io_outputWord[2];
  assign _T_248 = inner_io_outputWord[1];
  assign _T_249 = inner_io_outputWord[0];
  assign _T_251 = outputPieceBits == 6'h20;
  assign _T_254 = outputPieceBits + 6'h8;
  assign _T_255 = _T_254[5:0];
  assign _T_256 = _T_251 ? 6'h8 : _T_255;
  assign _T_260 = outputWriteAddr + 5'h1;
  assign _T_261 = _T_260[4:0];
  assign _T_262 = _T_251 ? _T_261 : outputWriteAddr;
  assign _T_264 = outputBits + 11'h8;
  assign _T_265 = _T_264[10:0];
  assign _GEN_63 = inner_io_outputValid ? _T_265 : outputBits;
  assign _GEN_64 = _T_241 ? _T_242 : outputMemBlock_31;
  assign _GEN_65 = _T_241 ? _T_243 : outputMemBlock_30;
  assign _GEN_66 = _T_241 ? _T_244 : outputMemBlock_29;
  assign _GEN_67 = _T_241 ? _T_245 : outputMemBlock_28;
  assign _GEN_68 = _T_241 ? _T_246 : outputMemBlock_27;
  assign _GEN_69 = _T_241 ? _T_247 : outputMemBlock_26;
  assign _GEN_70 = _T_241 ? _T_248 : outputMemBlock_25;
  assign _GEN_71 = _T_241 ? _T_249 : outputMemBlock_24;
  assign _GEN_72 = _T_241 ? outputMemBlock_8 : outputMemBlock_0;
  assign _GEN_73 = _T_241 ? outputMemBlock_9 : outputMemBlock_1;
  assign _GEN_74 = _T_241 ? outputMemBlock_10 : outputMemBlock_2;
  assign _GEN_75 = _T_241 ? outputMemBlock_11 : outputMemBlock_3;
  assign _GEN_76 = _T_241 ? outputMemBlock_12 : outputMemBlock_4;
  assign _GEN_77 = _T_241 ? outputMemBlock_13 : outputMemBlock_5;
  assign _GEN_78 = _T_241 ? outputMemBlock_14 : outputMemBlock_6;
  assign _GEN_79 = _T_241 ? outputMemBlock_15 : outputMemBlock_7;
  assign _GEN_80 = _T_241 ? outputMemBlock_16 : outputMemBlock_8;
  assign _GEN_81 = _T_241 ? outputMemBlock_17 : outputMemBlock_9;
  assign _GEN_82 = _T_241 ? outputMemBlock_18 : outputMemBlock_10;
  assign _GEN_83 = _T_241 ? outputMemBlock_19 : outputMemBlock_11;
  assign _GEN_84 = _T_241 ? outputMemBlock_20 : outputMemBlock_12;
  assign _GEN_85 = _T_241 ? outputMemBlock_21 : outputMemBlock_13;
  assign _GEN_86 = _T_241 ? outputMemBlock_22 : outputMemBlock_14;
  assign _GEN_87 = _T_241 ? outputMemBlock_23 : outputMemBlock_15;
  assign _GEN_88 = _T_241 ? outputMemBlock_24 : outputMemBlock_16;
  assign _GEN_89 = _T_241 ? outputMemBlock_25 : outputMemBlock_17;
  assign _GEN_90 = _T_241 ? outputMemBlock_26 : outputMemBlock_18;
  assign _GEN_91 = _T_241 ? outputMemBlock_27 : outputMemBlock_19;
  assign _GEN_92 = _T_241 ? outputMemBlock_28 : outputMemBlock_20;
  assign _GEN_93 = _T_241 ? outputMemBlock_29 : outputMemBlock_21;
  assign _GEN_94 = _T_241 ? outputMemBlock_30 : outputMemBlock_22;
  assign _GEN_95 = _T_241 ? outputMemBlock_31 : outputMemBlock_23;
  assign _GEN_96 = _T_241 ? _T_256 : outputPieceBits;
  assign _GEN_97 = _T_241 ? _T_262 : outputWriteAddr;
  assign _GEN_98 = _T_241 ? _GEN_63 : outputBits;
  assign _T_268 = {outputMemBlock_1,outputMemBlock_0};
  assign _T_269 = {outputMemBlock_3,outputMemBlock_2};
  assign _T_270 = {_T_269,_T_268};
  assign _T_271 = {outputMemBlock_5,outputMemBlock_4};
  assign _T_272 = {outputMemBlock_7,outputMemBlock_6};
  assign _T_273 = {_T_272,_T_271};
  assign _T_274 = {_T_273,_T_270};
  assign _T_275 = {outputMemBlock_9,outputMemBlock_8};
  assign _T_276 = {outputMemBlock_11,outputMemBlock_10};
  assign _T_277 = {_T_276,_T_275};
  assign _T_278 = {outputMemBlock_13,outputMemBlock_12};
  assign _T_279 = {outputMemBlock_15,outputMemBlock_14};
  assign _T_280 = {_T_279,_T_278};
  assign _T_281 = {_T_280,_T_277};
  assign _T_282 = {_T_281,_T_274};
  assign _T_283 = {outputMemBlock_17,outputMemBlock_16};
  assign _T_284 = {outputMemBlock_19,outputMemBlock_18};
  assign _T_285 = {_T_284,_T_283};
  assign _T_286 = {outputMemBlock_21,outputMemBlock_20};
  assign _T_287 = {outputMemBlock_23,outputMemBlock_22};
  assign _T_288 = {_T_287,_T_286};
  assign _T_289 = {_T_288,_T_285};
  assign _T_290 = {outputMemBlock_25,outputMemBlock_24};
  assign _T_291 = {outputMemBlock_27,outputMemBlock_26};
  assign _T_292 = {_T_291,_T_290};
  assign _T_293 = {outputMemBlock_29,outputMemBlock_28};
  assign _T_294 = {outputMemBlock_31,outputMemBlock_30};
  assign _T_295 = {_T_294,_T_293};
  assign _T_296 = {_T_295,_T_292};
  assign _T_297 = {_T_296,_T_289};
  assign _T_298 = {_T_297,_T_282};
  assign _T_305 = outputReadingStartedPrev == 1'h0;
  assign _T_309 = outputBits > 11'h0;
  assign _T_310 = inner_io_outputFinished & _T_309;
  assign _T_313 = _T_310 & _T_251;
  assign _T_314 = _T_231 | _T_313;
  assign _T_315 = _T_305 & _T_314;
  assign _GEN_99 = _T_315 ? 1'h1 : outputReadingStartedPrev;
  assign _T_318 = outputReadingStarted == 1'h0;
  assign _T_319 = outputReadingStartedPrev & _T_318;
  assign _GEN_100 = _T_319 ? 1'h1 : outputReadingStarted;
  assign _T_321 = io_outputMemBlockReady & outputReadingStarted;
  assign _T_323 = outputReadAddr == 5'h1f;
  assign _T_325 = _T_323 == 1'h0;
  assign _T_326 = _T_321 & _T_325;
  assign _T_328 = outputReadAddr + 5'h1;
  assign _T_329 = _T_328[4:0];
  assign _T_331 = outputReadAddr == 5'h0;
  assign _GEN_101 = _T_331 ? 11'h0 : _GEN_98;
  assign _GEN_102 = _T_326 ? _T_329 : outputReadAddr;
  assign _GEN_103 = _T_326 ? _GEN_101 : _GEN_98;
  assign _T_336 = outputBits == 11'h0;
  assign _T_337 = inner_io_outputFinished & _T_336;
  assign _T_340 = _T_337 & _T_331;
  assign _T_343 = outputReadingStarted & _T_323;
  assign _GEN_104 = _T_343 ? 1'h0 : _GEN_99;
  assign _GEN_105 = _T_343 ? 1'h0 : _GEN_100;
  assign _GEN_106 = _T_343 ? 5'h0 : _GEN_102;
  assign io_inputMemConsumed = _T_109;
  assign io_outputMemBlock = outputBram_io_b_dout;
  assign io_outputMemBlockValid = outputReadingStarted;
  assign io_outputBits = outputBits;
  assign io_outputFinished = _T_340;
  assign inner_io_inputWord = nextWord;
  assign inner_io_inputValid = _T_226;
  assign inner_io_inputFinished = _T_229;
  assign inner_io_outputReady = _T_233;
  assign inner_clock = clock;
  assign inner_reset = reset;
  assign inputBram_io_a_addr = io_inputMemIdx;
  assign inputBram_io_a_din = io_inputMemBlock;
  assign inputBram_io_a_wr = io_inputMemBlockValid;
  assign inputBram_io_b_addr = inputReadAddrFinal;
  assign inputBram_clock = clock;
  assign outputBram_io_a_addr = outputWriteAddr;
  assign outputBram_io_a_din = _T_298;
  assign outputBram_io_a_wr = _T_251;
  assign outputBram_io_b_addr = outputReadAddr;
  assign outputBram_clock = clock;
  assign inputReadAddrFinal = _GEN_4;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  inputMemBlock_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  inputMemBlock_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputMemBlock_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  inputMemBlock_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  inputMemBlock_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  inputMemBlock_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  inputMemBlock_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  inputMemBlock_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  inputMemBlock_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  inputMemBlock_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  inputMemBlock_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  inputMemBlock_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  inputMemBlock_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  inputMemBlock_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  inputMemBlock_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  inputMemBlock_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  inputMemBlock_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  inputMemBlock_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  inputMemBlock_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  inputMemBlock_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  inputMemBlock_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  inputMemBlock_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  inputMemBlock_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  inputMemBlock_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  inputMemBlock_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  inputMemBlock_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  inputMemBlock_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  inputMemBlock_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  inputMemBlock_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  inputMemBlock_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  inputMemBlock_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  inputMemBlock_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  inputPieceBitsRemaining = _RAND_32[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  inputBitsRemaining = _RAND_33[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  outputMemBlock_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  outputMemBlock_1 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  outputMemBlock_2 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  outputMemBlock_3 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  outputMemBlock_4 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  outputMemBlock_5 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  outputMemBlock_6 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  outputMemBlock_7 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  outputMemBlock_8 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  outputMemBlock_9 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  outputMemBlock_10 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  outputMemBlock_11 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  outputMemBlock_12 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  outputMemBlock_13 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  outputMemBlock_14 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  outputMemBlock_15 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  outputMemBlock_16 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  outputMemBlock_17 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  outputMemBlock_18 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  outputMemBlock_19 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  outputMemBlock_20 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  outputMemBlock_21 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  outputMemBlock_22 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  outputMemBlock_23 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  outputMemBlock_24 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  outputMemBlock_25 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  outputMemBlock_26 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  outputMemBlock_27 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  outputMemBlock_28 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  outputMemBlock_29 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  outputMemBlock_30 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  outputMemBlock_31 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  outputBits = _RAND_66[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  outputPieceBits = _RAND_67[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  inputReadAddr = _RAND_68[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  outputWriteAddr = _RAND_69[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  outputReadAddr = _RAND_70[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  outputReadingStartedPrev = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  outputReadingStarted = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_183) begin
      inputMemBlock_0 <= inputMemBlock_8;
    end else begin
      if (_T_121) begin
        inputMemBlock_0 <= _T_142;
      end
    end
    if (_T_183) begin
      inputMemBlock_1 <= inputMemBlock_9;
    end else begin
      if (_T_121) begin
        inputMemBlock_1 <= _T_143;
      end
    end
    if (_T_183) begin
      inputMemBlock_2 <= inputMemBlock_10;
    end else begin
      if (_T_121) begin
        inputMemBlock_2 <= _T_144;
      end
    end
    if (_T_183) begin
      inputMemBlock_3 <= inputMemBlock_11;
    end else begin
      if (_T_121) begin
        inputMemBlock_3 <= _T_145;
      end
    end
    if (_T_183) begin
      inputMemBlock_4 <= inputMemBlock_12;
    end else begin
      if (_T_121) begin
        inputMemBlock_4 <= _T_146;
      end
    end
    if (_T_183) begin
      inputMemBlock_5 <= inputMemBlock_13;
    end else begin
      if (_T_121) begin
        inputMemBlock_5 <= _T_147;
      end
    end
    if (_T_183) begin
      inputMemBlock_6 <= inputMemBlock_14;
    end else begin
      if (_T_121) begin
        inputMemBlock_6 <= _T_148;
      end
    end
    if (_T_183) begin
      inputMemBlock_7 <= inputMemBlock_15;
    end else begin
      if (_T_121) begin
        inputMemBlock_7 <= _T_149;
      end
    end
    if (_T_183) begin
      inputMemBlock_8 <= inputMemBlock_16;
    end else begin
      if (_T_121) begin
        inputMemBlock_8 <= _T_150;
      end
    end
    if (_T_183) begin
      inputMemBlock_9 <= inputMemBlock_17;
    end else begin
      if (_T_121) begin
        inputMemBlock_9 <= _T_151;
      end
    end
    if (_T_183) begin
      inputMemBlock_10 <= inputMemBlock_18;
    end else begin
      if (_T_121) begin
        inputMemBlock_10 <= _T_152;
      end
    end
    if (_T_183) begin
      inputMemBlock_11 <= inputMemBlock_19;
    end else begin
      if (_T_121) begin
        inputMemBlock_11 <= _T_153;
      end
    end
    if (_T_183) begin
      inputMemBlock_12 <= inputMemBlock_20;
    end else begin
      if (_T_121) begin
        inputMemBlock_12 <= _T_154;
      end
    end
    if (_T_183) begin
      inputMemBlock_13 <= inputMemBlock_21;
    end else begin
      if (_T_121) begin
        inputMemBlock_13 <= _T_155;
      end
    end
    if (_T_183) begin
      inputMemBlock_14 <= inputMemBlock_22;
    end else begin
      if (_T_121) begin
        inputMemBlock_14 <= _T_156;
      end
    end
    if (_T_183) begin
      inputMemBlock_15 <= inputMemBlock_23;
    end else begin
      if (_T_121) begin
        inputMemBlock_15 <= _T_157;
      end
    end
    if (_T_183) begin
      inputMemBlock_16 <= inputMemBlock_24;
    end else begin
      if (_T_121) begin
        inputMemBlock_16 <= _T_158;
      end
    end
    if (_T_183) begin
      inputMemBlock_17 <= inputMemBlock_25;
    end else begin
      if (_T_121) begin
        inputMemBlock_17 <= _T_159;
      end
    end
    if (_T_183) begin
      inputMemBlock_18 <= inputMemBlock_26;
    end else begin
      if (_T_121) begin
        inputMemBlock_18 <= _T_160;
      end
    end
    if (_T_183) begin
      inputMemBlock_19 <= inputMemBlock_27;
    end else begin
      if (_T_121) begin
        inputMemBlock_19 <= _T_161;
      end
    end
    if (_T_183) begin
      inputMemBlock_20 <= inputMemBlock_28;
    end else begin
      if (_T_121) begin
        inputMemBlock_20 <= _T_162;
      end
    end
    if (_T_183) begin
      inputMemBlock_21 <= inputMemBlock_29;
    end else begin
      if (_T_121) begin
        inputMemBlock_21 <= _T_163;
      end
    end
    if (_T_183) begin
      inputMemBlock_22 <= inputMemBlock_30;
    end else begin
      if (_T_121) begin
        inputMemBlock_22 <= _T_164;
      end
    end
    if (_T_183) begin
      inputMemBlock_23 <= inputMemBlock_31;
    end else begin
      if (_T_121) begin
        inputMemBlock_23 <= _T_165;
      end
    end
    if (_T_121) begin
      inputMemBlock_24 <= _T_166;
    end
    if (_T_121) begin
      inputMemBlock_25 <= _T_167;
    end
    if (_T_121) begin
      inputMemBlock_26 <= _T_168;
    end
    if (_T_121) begin
      inputMemBlock_27 <= _T_169;
    end
    if (_T_121) begin
      inputMemBlock_28 <= _T_170;
    end
    if (_T_121) begin
      inputMemBlock_29 <= _T_171;
    end
    if (_T_121) begin
      inputMemBlock_30 <= _T_172;
    end
    if (_T_121) begin
      inputMemBlock_31 <= _T_173;
    end
    if (reset) begin
      inputPieceBitsRemaining <= 6'h0;
    end else begin
      inputPieceBitsRemaining <= _GEN_37[5:0];
    end
    if (reset) begin
      inputBitsRemaining <= 11'h0;
    end else begin
      if (_T_183) begin
        inputBitsRemaining <= _T_127;
      end else begin
        if (_T_121) begin
          if (!(_T_107)) begin
            inputBitsRemaining <= _T_127;
          end
        end else begin
          if (_T_103) begin
            inputBitsRemaining <= io_inputBits;
          end
        end
      end
    end
    if (_T_241) begin
      outputMemBlock_0 <= outputMemBlock_8;
    end
    if (_T_241) begin
      outputMemBlock_1 <= outputMemBlock_9;
    end
    if (_T_241) begin
      outputMemBlock_2 <= outputMemBlock_10;
    end
    if (_T_241) begin
      outputMemBlock_3 <= outputMemBlock_11;
    end
    if (_T_241) begin
      outputMemBlock_4 <= outputMemBlock_12;
    end
    if (_T_241) begin
      outputMemBlock_5 <= outputMemBlock_13;
    end
    if (_T_241) begin
      outputMemBlock_6 <= outputMemBlock_14;
    end
    if (_T_241) begin
      outputMemBlock_7 <= outputMemBlock_15;
    end
    if (_T_241) begin
      outputMemBlock_8 <= outputMemBlock_16;
    end
    if (_T_241) begin
      outputMemBlock_9 <= outputMemBlock_17;
    end
    if (_T_241) begin
      outputMemBlock_10 <= outputMemBlock_18;
    end
    if (_T_241) begin
      outputMemBlock_11 <= outputMemBlock_19;
    end
    if (_T_241) begin
      outputMemBlock_12 <= outputMemBlock_20;
    end
    if (_T_241) begin
      outputMemBlock_13 <= outputMemBlock_21;
    end
    if (_T_241) begin
      outputMemBlock_14 <= outputMemBlock_22;
    end
    if (_T_241) begin
      outputMemBlock_15 <= outputMemBlock_23;
    end
    if (_T_241) begin
      outputMemBlock_16 <= outputMemBlock_24;
    end
    if (_T_241) begin
      outputMemBlock_17 <= outputMemBlock_25;
    end
    if (_T_241) begin
      outputMemBlock_18 <= outputMemBlock_26;
    end
    if (_T_241) begin
      outputMemBlock_19 <= outputMemBlock_27;
    end
    if (_T_241) begin
      outputMemBlock_20 <= outputMemBlock_28;
    end
    if (_T_241) begin
      outputMemBlock_21 <= outputMemBlock_29;
    end
    if (_T_241) begin
      outputMemBlock_22 <= outputMemBlock_30;
    end
    if (_T_241) begin
      outputMemBlock_23 <= outputMemBlock_31;
    end
    if (_T_241) begin
      outputMemBlock_24 <= _T_249;
    end
    if (_T_241) begin
      outputMemBlock_25 <= _T_248;
    end
    if (_T_241) begin
      outputMemBlock_26 <= _T_247;
    end
    if (_T_241) begin
      outputMemBlock_27 <= _T_246;
    end
    if (_T_241) begin
      outputMemBlock_28 <= _T_245;
    end
    if (_T_241) begin
      outputMemBlock_29 <= _T_244;
    end
    if (_T_241) begin
      outputMemBlock_30 <= _T_243;
    end
    if (_T_241) begin
      outputMemBlock_31 <= _T_242;
    end
    if (reset) begin
      outputBits <= 11'h0;
    end else begin
      if (_T_326) begin
        if (_T_331) begin
          outputBits <= 11'h0;
        end else begin
          if (_T_241) begin
            if (inner_io_outputValid) begin
              outputBits <= _T_265;
            end
          end
        end
      end else begin
        if (_T_241) begin
          if (inner_io_outputValid) begin
            outputBits <= _T_265;
          end
        end
      end
    end
    if (reset) begin
      outputPieceBits <= 6'h0;
    end else begin
      if (_T_241) begin
        if (_T_251) begin
          outputPieceBits <= 6'h8;
        end else begin
          outputPieceBits <= _T_255;
        end
      end
    end
    if (reset) begin
      inputReadAddr <= 5'h0;
    end else begin
      if (_T_121) begin
        if (!(_T_134)) begin
          inputReadAddr <= _T_137;
        end
      end
    end
    if (reset) begin
      outputWriteAddr <= 5'h0;
    end else begin
      if (_T_241) begin
        if (_T_251) begin
          outputWriteAddr <= _T_261;
        end
      end
    end
    if (reset) begin
      outputReadAddr <= 5'h0;
    end else begin
      if (_T_343) begin
        outputReadAddr <= 5'h0;
      end else begin
        if (_T_326) begin
          outputReadAddr <= _T_329;
        end
      end
    end
    if (reset) begin
      outputReadingStartedPrev <= 1'h0;
    end else begin
      if (_T_343) begin
        outputReadingStartedPrev <= 1'h0;
      end else begin
        if (_T_315) begin
          outputReadingStartedPrev <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputReadingStarted <= 1'h0;
    end else begin
      if (_T_343) begin
        outputReadingStarted <= 1'h0;
      end else begin
        if (_T_319) begin
          outputReadingStarted <= 1'h1;
        end
      end
    end
  end
endmodule
module StreamingCore(
  input         clock,
  input         reset,
  input  [31:0] io_metadataPtr,
  output [31:0] io_inputMemAddr,
  output        io_inputMemAddrValid,
  output        io_inputMemAddrsFinished,
  input  [31:0] io_inputMemBlock,
  input  [4:0]  io_inputMemIdx,
  input         io_inputMemBlockValid,
  output [31:0] io_outputMemAddr,
  output        io_outputMemAddrValid,
  input         io_outputMemAddrReady,
  output [31:0] io_outputMemBlock,
  output [4:0]  io_outputMemIdx,
  output        io_outputMemBlockValid,
  output        io_outputFinished
);
  wire  core_clock;
  wire  core_reset;
  wire [31:0] core_io_inputMemBlock;
  wire [4:0] core_io_inputMemIdx;
  wire  core_io_inputMemBlockValid;
  wire [10:0] core_io_inputBits;
  wire  core_io_inputMemConsumed;
  wire  core_io_inputFinished;
  wire [31:0] core_io_outputMemBlock;
  wire  core_io_outputMemBlockValid;
  wire  core_io_outputMemBlockReady;
  wire [10:0] core_io_outputBits;
  wire  core_io_outputFinished;
  reg  isInit;
  reg [31:0] _RAND_0;
  reg  initDone;
  reg [31:0] _RAND_1;
  reg [31:0] inputBitsRemaining;
  reg [31:0] _RAND_2;
  reg [31:0] outputBits;
  reg [31:0] _RAND_3;
  reg [4:0] outputBlockCounter;
  reg [31:0] _RAND_4;
  reg  outputLengthSent;
  reg [31:0] _RAND_5;
  reg [31:0] inputMemAddr;
  reg [31:0] _RAND_6;
  reg [31:0] outputMemAddr;
  reg [31:0] _RAND_7;
  reg [31:0] outputLenAddr;
  reg [31:0] _RAND_8;
  wire  _T_35;
  wire  _T_37;
  wire  _T_39;
  wire  _T_40;
  wire  _T_41;
  wire  _T_44;
  wire  _T_46;
  wire [31:0] _T_48;
  wire  _T_50;
  wire [31:0] _GEN_0;
  wire  _T_53;
  wire [31:0] _GEN_1;
  wire  _T_56;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_3;
  wire  _T_60;
  wire [32:0] _T_64;
  wire [31:0] _T_65;
  wire  _GEN_4;
  wire  _GEN_5;
  wire [31:0] _GEN_6;
  wire  _T_67;
  wire [32:0] _T_71;
  wire [32:0] _T_72;
  wire [31:0] _T_73;
  wire [31:0] _T_75;
  wire [32:0] _T_77;
  wire [31:0] _T_78;
  wire [31:0] _GEN_7;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [31:0] _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire [31:0] _GEN_15;
  wire [31:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [31:0] _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _T_81;
  reg  outputAddressAccepted;
  reg [31:0] _RAND_9;
  reg  outputAddressAcceptedNext;
  reg [31:0] _RAND_10;
  wire  _GEN_21;
  wire [31:0] _T_87;
  wire  _T_89;
  wire  _T_91;
  wire  _T_92;
  wire  _T_93;
  wire  _T_94;
  wire  _T_95;
  wire  _T_98;
  wire [31:0] _GEN_33;
  wire [32:0] _T_99;
  wire [31:0] _T_100;
  wire [31:0] _GEN_22;
  wire [31:0] _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire  _GEN_28;
  wire  _T_106;
  wire [5:0] _T_109;
  wire [4:0] _T_110;
  wire [4:0] _GEN_29;
  wire [4:0] _GEN_30;
  wire [31:0] outputBitsBlock;
  wire  _T_113;
  wire [31:0] tmp;
  wire [31:0] _T_116;
  wire  _T_119;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _T_124;
  InnerCore core (
    .clock(core_clock),
    .reset(core_reset),
    .io_inputMemBlock(core_io_inputMemBlock),
    .io_inputMemIdx(core_io_inputMemIdx),
    .io_inputMemBlockValid(core_io_inputMemBlockValid),
    .io_inputBits(core_io_inputBits),
    .io_inputMemConsumed(core_io_inputMemConsumed),
    .io_inputFinished(core_io_inputFinished),
    .io_outputMemBlock(core_io_outputMemBlock),
    .io_outputMemBlockValid(core_io_outputMemBlockValid),
    .io_outputMemBlockReady(core_io_outputMemBlockReady),
    .io_outputBits(core_io_outputBits),
    .io_outputFinished(core_io_outputFinished)
  );
  assign _T_35 = initDone & core_io_inputMemConsumed;
  assign _T_37 = inputBitsRemaining == 32'h0;
  assign _T_39 = _T_37 == 1'h0;
  assign _T_40 = _T_35 & _T_39;
  assign _T_41 = isInit | _T_40;
  assign _T_44 = io_inputMemBlockValid & initDone;
  assign _T_46 = inputBitsRemaining > 32'h400;
  assign _T_48 = _T_46 ? 32'h400 : inputBitsRemaining;
  assign _T_50 = io_inputMemIdx == 5'h0;
  assign _GEN_0 = _T_50 ? io_inputMemBlock : inputMemAddr;
  assign _T_53 = io_inputMemIdx == 5'h2;
  assign _GEN_1 = _T_53 ? io_inputMemBlock : inputBitsRemaining;
  assign _T_56 = io_inputMemIdx == 5'h4;
  assign _GEN_2 = _T_56 ? io_inputMemBlock : outputMemAddr;
  assign _GEN_3 = _T_56 ? io_inputMemBlock : outputLenAddr;
  assign _T_60 = io_inputMemIdx == 5'h1f;
  assign _T_64 = outputMemAddr + 32'h80;
  assign _T_65 = _T_64[31:0];
  assign _GEN_4 = _T_60 ? 1'h0 : isInit;
  assign _GEN_5 = _T_60 ? 1'h1 : initDone;
  assign _GEN_6 = _T_60 ? _T_65 : _GEN_2;
  assign _T_67 = io_inputMemIdx == 5'h1;
  assign _T_71 = inputBitsRemaining - 32'h400;
  assign _T_72 = $unsigned(_T_71);
  assign _T_73 = _T_72[31:0];
  assign _T_75 = _T_46 ? _T_73 : 32'h0;
  assign _T_77 = inputMemAddr + 32'h80;
  assign _T_78 = _T_77[31:0];
  assign _GEN_7 = _T_67 ? _T_75 : inputBitsRemaining;
  assign _GEN_8 = _T_67 ? _T_78 : inputMemAddr;
  assign _GEN_9 = isInit ? _GEN_0 : _GEN_8;
  assign _GEN_10 = isInit ? _GEN_1 : _GEN_7;
  assign _GEN_11 = isInit ? _GEN_6 : outputMemAddr;
  assign _GEN_12 = isInit ? _GEN_3 : outputLenAddr;
  assign _GEN_13 = isInit ? _GEN_4 : isInit;
  assign _GEN_14 = isInit ? _GEN_5 : initDone;
  assign _GEN_15 = io_inputMemBlockValid ? _GEN_9 : inputMemAddr;
  assign _GEN_16 = io_inputMemBlockValid ? _GEN_10 : inputBitsRemaining;
  assign _GEN_17 = io_inputMemBlockValid ? _GEN_11 : outputMemAddr;
  assign _GEN_18 = io_inputMemBlockValid ? _GEN_12 : outputLenAddr;
  assign _GEN_19 = io_inputMemBlockValid ? _GEN_13 : isInit;
  assign _GEN_20 = io_inputMemBlockValid ? _GEN_14 : initDone;
  assign _T_81 = initDone & _T_37;
  assign _GEN_21 = outputAddressAccepted ? 1'h1 : outputAddressAcceptedNext;
  assign _T_87 = core_io_outputFinished ? outputLenAddr : outputMemAddr;
  assign _T_89 = outputAddressAccepted == 1'h0;
  assign _T_91 = outputLengthSent == 1'h0;
  assign _T_92 = core_io_outputFinished & _T_91;
  assign _T_93 = core_io_outputMemBlockValid | _T_92;
  assign _T_94 = _T_89 & _T_93;
  assign _T_95 = io_outputMemAddrValid & io_outputMemAddrReady;
  assign _T_98 = core_io_outputFinished == 1'h0;
  assign _GEN_33 = {{21'd0}, core_io_outputBits};
  assign _T_99 = outputBits + _GEN_33;
  assign _T_100 = _T_99[31:0];
  assign _GEN_22 = _T_98 ? _T_100 : outputBits;
  assign _GEN_23 = _T_98 ? _T_65 : _GEN_17;
  assign _GEN_24 = _T_98 ? outputLengthSent : 1'h1;
  assign _GEN_25 = _T_95 ? 1'h1 : outputAddressAccepted;
  assign _GEN_26 = _T_95 ? _GEN_22 : outputBits;
  assign _GEN_27 = _T_95 ? _GEN_23 : _GEN_17;
  assign _GEN_28 = _T_95 ? _GEN_24 : outputLengthSent;
  assign _T_106 = outputBlockCounter == 5'h1f;
  assign _T_109 = outputBlockCounter + 5'h1;
  assign _T_110 = _T_109[4:0];
  assign _GEN_29 = _T_106 ? 5'h0 : _T_110;
  assign _GEN_30 = outputAddressAcceptedNext ? _GEN_29 : outputBlockCounter;
  assign _T_113 = outputBlockCounter == 5'h0;
  assign tmp = _T_113 ? outputBits : 32'h0;
  assign _T_116 = outputLengthSent ? outputBitsBlock : core_io_outputMemBlock;
  assign _T_119 = outputAddressAcceptedNext & _T_106;
  assign _GEN_31 = _T_119 ? 1'h0 : _GEN_25;
  assign _GEN_32 = _T_119 ? 1'h0 : _GEN_21;
  assign _T_124 = outputLengthSent & _T_89;
  assign io_inputMemAddr = inputMemAddr;
  assign io_inputMemAddrValid = _T_41;
  assign io_inputMemAddrsFinished = _T_37;
  assign io_outputMemAddr = _T_87;
  assign io_outputMemAddrValid = _T_94;
  assign io_outputMemBlock = _T_116;
  assign io_outputMemIdx = outputBlockCounter;
  assign io_outputMemBlockValid = outputAddressAcceptedNext;
  assign io_outputFinished = _T_124;
  assign core_io_inputMemBlock = io_inputMemBlock;
  assign core_io_inputMemIdx = io_inputMemIdx;
  assign core_io_inputMemBlockValid = _T_44;
  assign core_io_inputBits = _T_48[10:0];
  assign core_io_inputFinished = _T_81;
  assign core_io_outputMemBlockReady = outputAddressAccepted;
  assign core_clock = clock;
  assign core_reset = reset;
  assign outputBitsBlock = tmp;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  isInit = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  initDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  inputBitsRemaining = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  outputBits = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  outputBlockCounter = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputLengthSent = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  inputMemAddr = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  outputMemAddr = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  outputLenAddr = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  outputAddressAccepted = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  outputAddressAcceptedNext = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      isInit <= 1'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_60) begin
            isInit <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      initDone <= 1'h0;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_60) begin
            initDone <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBitsRemaining <= 32'h1;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_53) begin
            inputBitsRemaining <= io_inputMemBlock;
          end
        end else begin
          if (_T_67) begin
            if (_T_46) begin
              inputBitsRemaining <= _T_73;
            end else begin
              inputBitsRemaining <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      outputBits <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_98) begin
          outputBits <= _T_100;
        end
      end
    end
    if (reset) begin
      outputBlockCounter <= 5'h0;
    end else begin
      if (outputAddressAcceptedNext) begin
        if (_T_106) begin
          outputBlockCounter <= 5'h0;
        end else begin
          outputBlockCounter <= _T_110;
        end
      end
    end
    if (reset) begin
      outputLengthSent <= 1'h0;
    end else begin
      if (_T_95) begin
        if (!(_T_98)) begin
          outputLengthSent <= 1'h1;
        end
      end
    end
    if (reset) begin
      inputMemAddr <= io_metadataPtr;
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_50) begin
            inputMemAddr <= io_inputMemBlock;
          end
        end else begin
          if (_T_67) begin
            inputMemAddr <= _T_78;
          end
        end
      end
    end
    if (_T_95) begin
      if (_T_98) begin
        outputMemAddr <= _T_65;
      end else begin
        if (io_inputMemBlockValid) begin
          if (isInit) begin
            if (_T_60) begin
              outputMemAddr <= _T_65;
            end else begin
              if (_T_56) begin
                outputMemAddr <= io_inputMemBlock;
              end
            end
          end
        end
      end
    end else begin
      if (io_inputMemBlockValid) begin
        if (isInit) begin
          if (_T_60) begin
            outputMemAddr <= _T_65;
          end else begin
            if (_T_56) begin
              outputMemAddr <= io_inputMemBlock;
            end
          end
        end
      end
    end
    if (io_inputMemBlockValid) begin
      if (isInit) begin
        if (_T_56) begin
          outputLenAddr <= io_inputMemBlock;
        end
      end
    end
    if (reset) begin
      outputAddressAccepted <= 1'h0;
    end else begin
      if (_T_119) begin
        outputAddressAccepted <= 1'h0;
      end else begin
        if (_T_95) begin
          outputAddressAccepted <= 1'h1;
        end
      end
    end
    if (reset) begin
      outputAddressAcceptedNext <= 1'h0;
    end else begin
      if (_T_119) begin
        outputAddressAcceptedNext <= 1'h0;
      end else begin
        if (outputAddressAccepted) begin
          outputAddressAcceptedNext <= 1'h1;
        end
      end
    end
  end
endmodule
module StreamingWrapper(
  input          clock,
  input          reset,
  output [63:0]  io_inputMemAddrs_0,
  output [63:0]  io_inputMemAddrs_1,
  output [63:0]  io_inputMemAddrs_2,
  output [63:0]  io_inputMemAddrs_3,
  output         io_inputMemAddrValids_0,
  output         io_inputMemAddrValids_1,
  output         io_inputMemAddrValids_2,
  output         io_inputMemAddrValids_3,
  output [7:0]   io_inputMemAddrLens_0,
  output [7:0]   io_inputMemAddrLens_1,
  output [7:0]   io_inputMemAddrLens_2,
  output [7:0]   io_inputMemAddrLens_3,
  input          io_inputMemAddrReadys_0,
  input          io_inputMemAddrReadys_1,
  input          io_inputMemAddrReadys_2,
  input          io_inputMemAddrReadys_3,
  input  [511:0] io_inputMemBlocks_0,
  input  [511:0] io_inputMemBlocks_1,
  input  [511:0] io_inputMemBlocks_2,
  input  [511:0] io_inputMemBlocks_3,
  input          io_inputMemBlockValids_0,
  input          io_inputMemBlockValids_1,
  input          io_inputMemBlockValids_2,
  input          io_inputMemBlockValids_3,
  output         io_inputMemBlockReadys_0,
  output         io_inputMemBlockReadys_1,
  output         io_inputMemBlockReadys_2,
  output         io_inputMemBlockReadys_3,
  output [63:0]  io_outputMemAddrs_0,
  output [63:0]  io_outputMemAddrs_1,
  output [63:0]  io_outputMemAddrs_2,
  output [63:0]  io_outputMemAddrs_3,
  output         io_outputMemAddrValids_0,
  output         io_outputMemAddrValids_1,
  output         io_outputMemAddrValids_2,
  output         io_outputMemAddrValids_3,
  output [7:0]   io_outputMemAddrLens_0,
  output [7:0]   io_outputMemAddrLens_1,
  output [7:0]   io_outputMemAddrLens_2,
  output [7:0]   io_outputMemAddrLens_3,
  output [15:0]  io_outputMemAddrIds_0,
  output [15:0]  io_outputMemAddrIds_1,
  output [15:0]  io_outputMemAddrIds_2,
  output [15:0]  io_outputMemAddrIds_3,
  input          io_outputMemAddrReadys_0,
  input          io_outputMemAddrReadys_1,
  input          io_outputMemAddrReadys_2,
  input          io_outputMemAddrReadys_3,
  output [511:0] io_outputMemBlocks_0,
  output [511:0] io_outputMemBlocks_1,
  output [511:0] io_outputMemBlocks_2,
  output [511:0] io_outputMemBlocks_3,
  output         io_outputMemBlockValids_0,
  output         io_outputMemBlockValids_1,
  output         io_outputMemBlockValids_2,
  output         io_outputMemBlockValids_3,
  output         io_outputMemBlockLasts_0,
  output         io_outputMemBlockLasts_1,
  output         io_outputMemBlockLasts_2,
  output         io_outputMemBlockLasts_3,
  input          io_outputMemBlockReadys_0,
  input          io_outputMemBlockReadys_1,
  input          io_outputMemBlockReadys_2,
  input          io_outputMemBlockReadys_3,
  output         io_finished
);
  wire  mc_clock;
  wire  mc_reset;
  wire [63:0] mc_io_axi_inputMemAddrs_0;
  wire [63:0] mc_io_axi_inputMemAddrs_1;
  wire [63:0] mc_io_axi_inputMemAddrs_2;
  wire [63:0] mc_io_axi_inputMemAddrs_3;
  wire  mc_io_axi_inputMemAddrValids_0;
  wire  mc_io_axi_inputMemAddrValids_1;
  wire  mc_io_axi_inputMemAddrValids_2;
  wire  mc_io_axi_inputMemAddrValids_3;
  wire [7:0] mc_io_axi_inputMemAddrLens_0;
  wire [7:0] mc_io_axi_inputMemAddrLens_1;
  wire [7:0] mc_io_axi_inputMemAddrLens_2;
  wire [7:0] mc_io_axi_inputMemAddrLens_3;
  wire  mc_io_axi_inputMemAddrReadys_0;
  wire  mc_io_axi_inputMemAddrReadys_1;
  wire  mc_io_axi_inputMemAddrReadys_2;
  wire  mc_io_axi_inputMemAddrReadys_3;
  wire [511:0] mc_io_axi_inputMemBlocks_0;
  wire [511:0] mc_io_axi_inputMemBlocks_1;
  wire [511:0] mc_io_axi_inputMemBlocks_2;
  wire [511:0] mc_io_axi_inputMemBlocks_3;
  wire  mc_io_axi_inputMemBlockValids_0;
  wire  mc_io_axi_inputMemBlockValids_1;
  wire  mc_io_axi_inputMemBlockValids_2;
  wire  mc_io_axi_inputMemBlockValids_3;
  wire  mc_io_axi_inputMemBlockReadys_0;
  wire  mc_io_axi_inputMemBlockReadys_1;
  wire  mc_io_axi_inputMemBlockReadys_2;
  wire  mc_io_axi_inputMemBlockReadys_3;
  wire [63:0] mc_io_axi_outputMemAddrs_0;
  wire [63:0] mc_io_axi_outputMemAddrs_1;
  wire [63:0] mc_io_axi_outputMemAddrs_2;
  wire [63:0] mc_io_axi_outputMemAddrs_3;
  wire  mc_io_axi_outputMemAddrValids_0;
  wire  mc_io_axi_outputMemAddrValids_1;
  wire  mc_io_axi_outputMemAddrValids_2;
  wire  mc_io_axi_outputMemAddrValids_3;
  wire [7:0] mc_io_axi_outputMemAddrLens_0;
  wire [7:0] mc_io_axi_outputMemAddrLens_1;
  wire [7:0] mc_io_axi_outputMemAddrLens_2;
  wire [7:0] mc_io_axi_outputMemAddrLens_3;
  wire [15:0] mc_io_axi_outputMemAddrIds_0;
  wire [15:0] mc_io_axi_outputMemAddrIds_1;
  wire [15:0] mc_io_axi_outputMemAddrIds_2;
  wire [15:0] mc_io_axi_outputMemAddrIds_3;
  wire  mc_io_axi_outputMemAddrReadys_0;
  wire  mc_io_axi_outputMemAddrReadys_1;
  wire  mc_io_axi_outputMemAddrReadys_2;
  wire  mc_io_axi_outputMemAddrReadys_3;
  wire [511:0] mc_io_axi_outputMemBlocks_0;
  wire [511:0] mc_io_axi_outputMemBlocks_1;
  wire [511:0] mc_io_axi_outputMemBlocks_2;
  wire [511:0] mc_io_axi_outputMemBlocks_3;
  wire  mc_io_axi_outputMemBlockValids_0;
  wire  mc_io_axi_outputMemBlockValids_1;
  wire  mc_io_axi_outputMemBlockValids_2;
  wire  mc_io_axi_outputMemBlockValids_3;
  wire  mc_io_axi_outputMemBlockLasts_0;
  wire  mc_io_axi_outputMemBlockLasts_1;
  wire  mc_io_axi_outputMemBlockLasts_2;
  wire  mc_io_axi_outputMemBlockLasts_3;
  wire  mc_io_axi_outputMemBlockReadys_0;
  wire  mc_io_axi_outputMemBlockReadys_1;
  wire  mc_io_axi_outputMemBlockReadys_2;
  wire  mc_io_axi_outputMemBlockReadys_3;
  wire  mc_io_axi_finished;
  wire [31:0] mc_io_streamingCores_0_metadataPtr;
  wire [31:0] mc_io_streamingCores_0_inputMemAddr;
  wire  mc_io_streamingCores_0_inputMemAddrValid;
  wire  mc_io_streamingCores_0_inputMemAddrsFinished;
  wire [31:0] mc_io_streamingCores_0_inputMemBlock;
  wire [4:0] mc_io_streamingCores_0_inputMemIdx;
  wire  mc_io_streamingCores_0_inputMemBlockValid;
  wire [31:0] mc_io_streamingCores_0_outputMemAddr;
  wire  mc_io_streamingCores_0_outputMemAddrValid;
  wire  mc_io_streamingCores_0_outputMemAddrReady;
  wire [31:0] mc_io_streamingCores_0_outputMemBlock;
  wire [4:0] mc_io_streamingCores_0_outputMemIdx;
  wire  mc_io_streamingCores_0_outputMemBlockValid;
  wire  mc_io_streamingCores_0_outputFinished;
  wire [31:0] mc_io_streamingCores_1_metadataPtr;
  wire [31:0] mc_io_streamingCores_1_inputMemAddr;
  wire  mc_io_streamingCores_1_inputMemAddrValid;
  wire  mc_io_streamingCores_1_inputMemAddrsFinished;
  wire [31:0] mc_io_streamingCores_1_inputMemBlock;
  wire [4:0] mc_io_streamingCores_1_inputMemIdx;
  wire  mc_io_streamingCores_1_inputMemBlockValid;
  wire [31:0] mc_io_streamingCores_1_outputMemAddr;
  wire  mc_io_streamingCores_1_outputMemAddrValid;
  wire  mc_io_streamingCores_1_outputMemAddrReady;
  wire [31:0] mc_io_streamingCores_1_outputMemBlock;
  wire [4:0] mc_io_streamingCores_1_outputMemIdx;
  wire  mc_io_streamingCores_1_outputMemBlockValid;
  wire  mc_io_streamingCores_1_outputFinished;
  wire [31:0] mc_io_streamingCores_2_metadataPtr;
  wire [31:0] mc_io_streamingCores_2_inputMemAddr;
  wire  mc_io_streamingCores_2_inputMemAddrValid;
  wire  mc_io_streamingCores_2_inputMemAddrsFinished;
  wire [31:0] mc_io_streamingCores_2_inputMemBlock;
  wire [4:0] mc_io_streamingCores_2_inputMemIdx;
  wire  mc_io_streamingCores_2_inputMemBlockValid;
  wire [31:0] mc_io_streamingCores_2_outputMemAddr;
  wire  mc_io_streamingCores_2_outputMemAddrValid;
  wire  mc_io_streamingCores_2_outputMemAddrReady;
  wire [31:0] mc_io_streamingCores_2_outputMemBlock;
  wire [4:0] mc_io_streamingCores_2_outputMemIdx;
  wire  mc_io_streamingCores_2_outputMemBlockValid;
  wire  mc_io_streamingCores_2_outputFinished;
  wire [31:0] mc_io_streamingCores_3_metadataPtr;
  wire [31:0] mc_io_streamingCores_3_inputMemAddr;
  wire  mc_io_streamingCores_3_inputMemAddrValid;
  wire  mc_io_streamingCores_3_inputMemAddrsFinished;
  wire [31:0] mc_io_streamingCores_3_inputMemBlock;
  wire [4:0] mc_io_streamingCores_3_inputMemIdx;
  wire  mc_io_streamingCores_3_inputMemBlockValid;
  wire [31:0] mc_io_streamingCores_3_outputMemAddr;
  wire  mc_io_streamingCores_3_outputMemAddrValid;
  wire  mc_io_streamingCores_3_outputMemAddrReady;
  wire [31:0] mc_io_streamingCores_3_outputMemBlock;
  wire [4:0] mc_io_streamingCores_3_outputMemIdx;
  wire  mc_io_streamingCores_3_outputMemBlockValid;
  wire  mc_io_streamingCores_3_outputFinished;
  wire  StreamingCore_clock;
  wire  StreamingCore_reset;
  wire [31:0] StreamingCore_io_metadataPtr;
  wire [31:0] StreamingCore_io_inputMemAddr;
  wire  StreamingCore_io_inputMemAddrValid;
  wire  StreamingCore_io_inputMemAddrsFinished;
  wire [31:0] StreamingCore_io_inputMemBlock;
  wire [4:0] StreamingCore_io_inputMemIdx;
  wire  StreamingCore_io_inputMemBlockValid;
  wire [31:0] StreamingCore_io_outputMemAddr;
  wire  StreamingCore_io_outputMemAddrValid;
  wire  StreamingCore_io_outputMemAddrReady;
  wire [31:0] StreamingCore_io_outputMemBlock;
  wire [4:0] StreamingCore_io_outputMemIdx;
  wire  StreamingCore_io_outputMemBlockValid;
  wire  StreamingCore_io_outputFinished;
  wire  StreamingCore_1_clock;
  wire  StreamingCore_1_reset;
  wire [31:0] StreamingCore_1_io_metadataPtr;
  wire [31:0] StreamingCore_1_io_inputMemAddr;
  wire  StreamingCore_1_io_inputMemAddrValid;
  wire  StreamingCore_1_io_inputMemAddrsFinished;
  wire [31:0] StreamingCore_1_io_inputMemBlock;
  wire [4:0] StreamingCore_1_io_inputMemIdx;
  wire  StreamingCore_1_io_inputMemBlockValid;
  wire [31:0] StreamingCore_1_io_outputMemAddr;
  wire  StreamingCore_1_io_outputMemAddrValid;
  wire  StreamingCore_1_io_outputMemAddrReady;
  wire [31:0] StreamingCore_1_io_outputMemBlock;
  wire [4:0] StreamingCore_1_io_outputMemIdx;
  wire  StreamingCore_1_io_outputMemBlockValid;
  wire  StreamingCore_1_io_outputFinished;
  wire  StreamingCore_2_clock;
  wire  StreamingCore_2_reset;
  wire [31:0] StreamingCore_2_io_metadataPtr;
  wire [31:0] StreamingCore_2_io_inputMemAddr;
  wire  StreamingCore_2_io_inputMemAddrValid;
  wire  StreamingCore_2_io_inputMemAddrsFinished;
  wire [31:0] StreamingCore_2_io_inputMemBlock;
  wire [4:0] StreamingCore_2_io_inputMemIdx;
  wire  StreamingCore_2_io_inputMemBlockValid;
  wire [31:0] StreamingCore_2_io_outputMemAddr;
  wire  StreamingCore_2_io_outputMemAddrValid;
  wire  StreamingCore_2_io_outputMemAddrReady;
  wire [31:0] StreamingCore_2_io_outputMemBlock;
  wire [4:0] StreamingCore_2_io_outputMemIdx;
  wire  StreamingCore_2_io_outputMemBlockValid;
  wire  StreamingCore_2_io_outputFinished;
  wire  StreamingCore_3_clock;
  wire  StreamingCore_3_reset;
  wire [31:0] StreamingCore_3_io_metadataPtr;
  wire [31:0] StreamingCore_3_io_inputMemAddr;
  wire  StreamingCore_3_io_inputMemAddrValid;
  wire  StreamingCore_3_io_inputMemAddrsFinished;
  wire [31:0] StreamingCore_3_io_inputMemBlock;
  wire [4:0] StreamingCore_3_io_inputMemIdx;
  wire  StreamingCore_3_io_inputMemBlockValid;
  wire [31:0] StreamingCore_3_io_outputMemAddr;
  wire  StreamingCore_3_io_outputMemAddrValid;
  wire  StreamingCore_3_io_outputMemAddrReady;
  wire [31:0] StreamingCore_3_io_outputMemBlock;
  wire [4:0] StreamingCore_3_io_outputMemIdx;
  wire  StreamingCore_3_io_outputMemBlockValid;
  wire  StreamingCore_3_io_outputFinished;
  StreamingMemoryController mc (
    .clock(mc_clock),
    .reset(mc_reset),
    .io_axi_inputMemAddrs_0(mc_io_axi_inputMemAddrs_0),
    .io_axi_inputMemAddrs_1(mc_io_axi_inputMemAddrs_1),
    .io_axi_inputMemAddrs_2(mc_io_axi_inputMemAddrs_2),
    .io_axi_inputMemAddrs_3(mc_io_axi_inputMemAddrs_3),
    .io_axi_inputMemAddrValids_0(mc_io_axi_inputMemAddrValids_0),
    .io_axi_inputMemAddrValids_1(mc_io_axi_inputMemAddrValids_1),
    .io_axi_inputMemAddrValids_2(mc_io_axi_inputMemAddrValids_2),
    .io_axi_inputMemAddrValids_3(mc_io_axi_inputMemAddrValids_3),
    .io_axi_inputMemAddrLens_0(mc_io_axi_inputMemAddrLens_0),
    .io_axi_inputMemAddrLens_1(mc_io_axi_inputMemAddrLens_1),
    .io_axi_inputMemAddrLens_2(mc_io_axi_inputMemAddrLens_2),
    .io_axi_inputMemAddrLens_3(mc_io_axi_inputMemAddrLens_3),
    .io_axi_inputMemAddrReadys_0(mc_io_axi_inputMemAddrReadys_0),
    .io_axi_inputMemAddrReadys_1(mc_io_axi_inputMemAddrReadys_1),
    .io_axi_inputMemAddrReadys_2(mc_io_axi_inputMemAddrReadys_2),
    .io_axi_inputMemAddrReadys_3(mc_io_axi_inputMemAddrReadys_3),
    .io_axi_inputMemBlocks_0(mc_io_axi_inputMemBlocks_0),
    .io_axi_inputMemBlocks_1(mc_io_axi_inputMemBlocks_1),
    .io_axi_inputMemBlocks_2(mc_io_axi_inputMemBlocks_2),
    .io_axi_inputMemBlocks_3(mc_io_axi_inputMemBlocks_3),
    .io_axi_inputMemBlockValids_0(mc_io_axi_inputMemBlockValids_0),
    .io_axi_inputMemBlockValids_1(mc_io_axi_inputMemBlockValids_1),
    .io_axi_inputMemBlockValids_2(mc_io_axi_inputMemBlockValids_2),
    .io_axi_inputMemBlockValids_3(mc_io_axi_inputMemBlockValids_3),
    .io_axi_inputMemBlockReadys_0(mc_io_axi_inputMemBlockReadys_0),
    .io_axi_inputMemBlockReadys_1(mc_io_axi_inputMemBlockReadys_1),
    .io_axi_inputMemBlockReadys_2(mc_io_axi_inputMemBlockReadys_2),
    .io_axi_inputMemBlockReadys_3(mc_io_axi_inputMemBlockReadys_3),
    .io_axi_outputMemAddrs_0(mc_io_axi_outputMemAddrs_0),
    .io_axi_outputMemAddrs_1(mc_io_axi_outputMemAddrs_1),
    .io_axi_outputMemAddrs_2(mc_io_axi_outputMemAddrs_2),
    .io_axi_outputMemAddrs_3(mc_io_axi_outputMemAddrs_3),
    .io_axi_outputMemAddrValids_0(mc_io_axi_outputMemAddrValids_0),
    .io_axi_outputMemAddrValids_1(mc_io_axi_outputMemAddrValids_1),
    .io_axi_outputMemAddrValids_2(mc_io_axi_outputMemAddrValids_2),
    .io_axi_outputMemAddrValids_3(mc_io_axi_outputMemAddrValids_3),
    .io_axi_outputMemAddrLens_0(mc_io_axi_outputMemAddrLens_0),
    .io_axi_outputMemAddrLens_1(mc_io_axi_outputMemAddrLens_1),
    .io_axi_outputMemAddrLens_2(mc_io_axi_outputMemAddrLens_2),
    .io_axi_outputMemAddrLens_3(mc_io_axi_outputMemAddrLens_3),
    .io_axi_outputMemAddrIds_0(mc_io_axi_outputMemAddrIds_0),
    .io_axi_outputMemAddrIds_1(mc_io_axi_outputMemAddrIds_1),
    .io_axi_outputMemAddrIds_2(mc_io_axi_outputMemAddrIds_2),
    .io_axi_outputMemAddrIds_3(mc_io_axi_outputMemAddrIds_3),
    .io_axi_outputMemAddrReadys_0(mc_io_axi_outputMemAddrReadys_0),
    .io_axi_outputMemAddrReadys_1(mc_io_axi_outputMemAddrReadys_1),
    .io_axi_outputMemAddrReadys_2(mc_io_axi_outputMemAddrReadys_2),
    .io_axi_outputMemAddrReadys_3(mc_io_axi_outputMemAddrReadys_3),
    .io_axi_outputMemBlocks_0(mc_io_axi_outputMemBlocks_0),
    .io_axi_outputMemBlocks_1(mc_io_axi_outputMemBlocks_1),
    .io_axi_outputMemBlocks_2(mc_io_axi_outputMemBlocks_2),
    .io_axi_outputMemBlocks_3(mc_io_axi_outputMemBlocks_3),
    .io_axi_outputMemBlockValids_0(mc_io_axi_outputMemBlockValids_0),
    .io_axi_outputMemBlockValids_1(mc_io_axi_outputMemBlockValids_1),
    .io_axi_outputMemBlockValids_2(mc_io_axi_outputMemBlockValids_2),
    .io_axi_outputMemBlockValids_3(mc_io_axi_outputMemBlockValids_3),
    .io_axi_outputMemBlockLasts_0(mc_io_axi_outputMemBlockLasts_0),
    .io_axi_outputMemBlockLasts_1(mc_io_axi_outputMemBlockLasts_1),
    .io_axi_outputMemBlockLasts_2(mc_io_axi_outputMemBlockLasts_2),
    .io_axi_outputMemBlockLasts_3(mc_io_axi_outputMemBlockLasts_3),
    .io_axi_outputMemBlockReadys_0(mc_io_axi_outputMemBlockReadys_0),
    .io_axi_outputMemBlockReadys_1(mc_io_axi_outputMemBlockReadys_1),
    .io_axi_outputMemBlockReadys_2(mc_io_axi_outputMemBlockReadys_2),
    .io_axi_outputMemBlockReadys_3(mc_io_axi_outputMemBlockReadys_3),
    .io_axi_finished(mc_io_axi_finished),
    .io_streamingCores_0_metadataPtr(mc_io_streamingCores_0_metadataPtr),
    .io_streamingCores_0_inputMemAddr(mc_io_streamingCores_0_inputMemAddr),
    .io_streamingCores_0_inputMemAddrValid(mc_io_streamingCores_0_inputMemAddrValid),
    .io_streamingCores_0_inputMemAddrsFinished(mc_io_streamingCores_0_inputMemAddrsFinished),
    .io_streamingCores_0_inputMemBlock(mc_io_streamingCores_0_inputMemBlock),
    .io_streamingCores_0_inputMemIdx(mc_io_streamingCores_0_inputMemIdx),
    .io_streamingCores_0_inputMemBlockValid(mc_io_streamingCores_0_inputMemBlockValid),
    .io_streamingCores_0_outputMemAddr(mc_io_streamingCores_0_outputMemAddr),
    .io_streamingCores_0_outputMemAddrValid(mc_io_streamingCores_0_outputMemAddrValid),
    .io_streamingCores_0_outputMemAddrReady(mc_io_streamingCores_0_outputMemAddrReady),
    .io_streamingCores_0_outputMemBlock(mc_io_streamingCores_0_outputMemBlock),
    .io_streamingCores_0_outputMemIdx(mc_io_streamingCores_0_outputMemIdx),
    .io_streamingCores_0_outputMemBlockValid(mc_io_streamingCores_0_outputMemBlockValid),
    .io_streamingCores_0_outputFinished(mc_io_streamingCores_0_outputFinished),
    .io_streamingCores_1_metadataPtr(mc_io_streamingCores_1_metadataPtr),
    .io_streamingCores_1_inputMemAddr(mc_io_streamingCores_1_inputMemAddr),
    .io_streamingCores_1_inputMemAddrValid(mc_io_streamingCores_1_inputMemAddrValid),
    .io_streamingCores_1_inputMemAddrsFinished(mc_io_streamingCores_1_inputMemAddrsFinished),
    .io_streamingCores_1_inputMemBlock(mc_io_streamingCores_1_inputMemBlock),
    .io_streamingCores_1_inputMemIdx(mc_io_streamingCores_1_inputMemIdx),
    .io_streamingCores_1_inputMemBlockValid(mc_io_streamingCores_1_inputMemBlockValid),
    .io_streamingCores_1_outputMemAddr(mc_io_streamingCores_1_outputMemAddr),
    .io_streamingCores_1_outputMemAddrValid(mc_io_streamingCores_1_outputMemAddrValid),
    .io_streamingCores_1_outputMemAddrReady(mc_io_streamingCores_1_outputMemAddrReady),
    .io_streamingCores_1_outputMemBlock(mc_io_streamingCores_1_outputMemBlock),
    .io_streamingCores_1_outputMemIdx(mc_io_streamingCores_1_outputMemIdx),
    .io_streamingCores_1_outputMemBlockValid(mc_io_streamingCores_1_outputMemBlockValid),
    .io_streamingCores_1_outputFinished(mc_io_streamingCores_1_outputFinished),
    .io_streamingCores_2_metadataPtr(mc_io_streamingCores_2_metadataPtr),
    .io_streamingCores_2_inputMemAddr(mc_io_streamingCores_2_inputMemAddr),
    .io_streamingCores_2_inputMemAddrValid(mc_io_streamingCores_2_inputMemAddrValid),
    .io_streamingCores_2_inputMemAddrsFinished(mc_io_streamingCores_2_inputMemAddrsFinished),
    .io_streamingCores_2_inputMemBlock(mc_io_streamingCores_2_inputMemBlock),
    .io_streamingCores_2_inputMemIdx(mc_io_streamingCores_2_inputMemIdx),
    .io_streamingCores_2_inputMemBlockValid(mc_io_streamingCores_2_inputMemBlockValid),
    .io_streamingCores_2_outputMemAddr(mc_io_streamingCores_2_outputMemAddr),
    .io_streamingCores_2_outputMemAddrValid(mc_io_streamingCores_2_outputMemAddrValid),
    .io_streamingCores_2_outputMemAddrReady(mc_io_streamingCores_2_outputMemAddrReady),
    .io_streamingCores_2_outputMemBlock(mc_io_streamingCores_2_outputMemBlock),
    .io_streamingCores_2_outputMemIdx(mc_io_streamingCores_2_outputMemIdx),
    .io_streamingCores_2_outputMemBlockValid(mc_io_streamingCores_2_outputMemBlockValid),
    .io_streamingCores_2_outputFinished(mc_io_streamingCores_2_outputFinished),
    .io_streamingCores_3_metadataPtr(mc_io_streamingCores_3_metadataPtr),
    .io_streamingCores_3_inputMemAddr(mc_io_streamingCores_3_inputMemAddr),
    .io_streamingCores_3_inputMemAddrValid(mc_io_streamingCores_3_inputMemAddrValid),
    .io_streamingCores_3_inputMemAddrsFinished(mc_io_streamingCores_3_inputMemAddrsFinished),
    .io_streamingCores_3_inputMemBlock(mc_io_streamingCores_3_inputMemBlock),
    .io_streamingCores_3_inputMemIdx(mc_io_streamingCores_3_inputMemIdx),
    .io_streamingCores_3_inputMemBlockValid(mc_io_streamingCores_3_inputMemBlockValid),
    .io_streamingCores_3_outputMemAddr(mc_io_streamingCores_3_outputMemAddr),
    .io_streamingCores_3_outputMemAddrValid(mc_io_streamingCores_3_outputMemAddrValid),
    .io_streamingCores_3_outputMemAddrReady(mc_io_streamingCores_3_outputMemAddrReady),
    .io_streamingCores_3_outputMemBlock(mc_io_streamingCores_3_outputMemBlock),
    .io_streamingCores_3_outputMemIdx(mc_io_streamingCores_3_outputMemIdx),
    .io_streamingCores_3_outputMemBlockValid(mc_io_streamingCores_3_outputMemBlockValid),
    .io_streamingCores_3_outputFinished(mc_io_streamingCores_3_outputFinished)
  );
  StreamingCore StreamingCore (
    .clock(StreamingCore_clock),
    .reset(StreamingCore_reset),
    .io_metadataPtr(StreamingCore_io_metadataPtr),
    .io_inputMemAddr(StreamingCore_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_io_inputMemAddrValid),
    .io_inputMemAddrsFinished(StreamingCore_io_inputMemAddrsFinished),
    .io_inputMemBlock(StreamingCore_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_io_inputMemBlockValid),
    .io_outputMemAddr(StreamingCore_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_io_outputMemBlockValid),
    .io_outputFinished(StreamingCore_io_outputFinished)
  );
  StreamingCore StreamingCore_1 (
    .clock(StreamingCore_1_clock),
    .reset(StreamingCore_1_reset),
    .io_metadataPtr(StreamingCore_1_io_metadataPtr),
    .io_inputMemAddr(StreamingCore_1_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_1_io_inputMemAddrValid),
    .io_inputMemAddrsFinished(StreamingCore_1_io_inputMemAddrsFinished),
    .io_inputMemBlock(StreamingCore_1_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_1_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_1_io_inputMemBlockValid),
    .io_outputMemAddr(StreamingCore_1_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_1_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_1_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_1_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_1_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_1_io_outputMemBlockValid),
    .io_outputFinished(StreamingCore_1_io_outputFinished)
  );
  StreamingCore StreamingCore_2 (
    .clock(StreamingCore_2_clock),
    .reset(StreamingCore_2_reset),
    .io_metadataPtr(StreamingCore_2_io_metadataPtr),
    .io_inputMemAddr(StreamingCore_2_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_2_io_inputMemAddrValid),
    .io_inputMemAddrsFinished(StreamingCore_2_io_inputMemAddrsFinished),
    .io_inputMemBlock(StreamingCore_2_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_2_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_2_io_inputMemBlockValid),
    .io_outputMemAddr(StreamingCore_2_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_2_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_2_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_2_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_2_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_2_io_outputMemBlockValid),
    .io_outputFinished(StreamingCore_2_io_outputFinished)
  );
  StreamingCore StreamingCore_3 (
    .clock(StreamingCore_3_clock),
    .reset(StreamingCore_3_reset),
    .io_metadataPtr(StreamingCore_3_io_metadataPtr),
    .io_inputMemAddr(StreamingCore_3_io_inputMemAddr),
    .io_inputMemAddrValid(StreamingCore_3_io_inputMemAddrValid),
    .io_inputMemAddrsFinished(StreamingCore_3_io_inputMemAddrsFinished),
    .io_inputMemBlock(StreamingCore_3_io_inputMemBlock),
    .io_inputMemIdx(StreamingCore_3_io_inputMemIdx),
    .io_inputMemBlockValid(StreamingCore_3_io_inputMemBlockValid),
    .io_outputMemAddr(StreamingCore_3_io_outputMemAddr),
    .io_outputMemAddrValid(StreamingCore_3_io_outputMemAddrValid),
    .io_outputMemAddrReady(StreamingCore_3_io_outputMemAddrReady),
    .io_outputMemBlock(StreamingCore_3_io_outputMemBlock),
    .io_outputMemIdx(StreamingCore_3_io_outputMemIdx),
    .io_outputMemBlockValid(StreamingCore_3_io_outputMemBlockValid),
    .io_outputFinished(StreamingCore_3_io_outputFinished)
  );
  assign io_inputMemAddrs_0 = mc_io_axi_inputMemAddrs_0;
  assign io_inputMemAddrs_1 = mc_io_axi_inputMemAddrs_1;
  assign io_inputMemAddrs_2 = mc_io_axi_inputMemAddrs_2;
  assign io_inputMemAddrs_3 = mc_io_axi_inputMemAddrs_3;
  assign io_inputMemAddrValids_0 = mc_io_axi_inputMemAddrValids_0;
  assign io_inputMemAddrValids_1 = mc_io_axi_inputMemAddrValids_1;
  assign io_inputMemAddrValids_2 = mc_io_axi_inputMemAddrValids_2;
  assign io_inputMemAddrValids_3 = mc_io_axi_inputMemAddrValids_3;
  assign io_inputMemAddrLens_0 = mc_io_axi_inputMemAddrLens_0;
  assign io_inputMemAddrLens_1 = mc_io_axi_inputMemAddrLens_1;
  assign io_inputMemAddrLens_2 = mc_io_axi_inputMemAddrLens_2;
  assign io_inputMemAddrLens_3 = mc_io_axi_inputMemAddrLens_3;
  assign io_inputMemBlockReadys_0 = mc_io_axi_inputMemBlockReadys_0;
  assign io_inputMemBlockReadys_1 = mc_io_axi_inputMemBlockReadys_1;
  assign io_inputMemBlockReadys_2 = mc_io_axi_inputMemBlockReadys_2;
  assign io_inputMemBlockReadys_3 = mc_io_axi_inputMemBlockReadys_3;
  assign io_outputMemAddrs_0 = mc_io_axi_outputMemAddrs_0;
  assign io_outputMemAddrs_1 = mc_io_axi_outputMemAddrs_1;
  assign io_outputMemAddrs_2 = mc_io_axi_outputMemAddrs_2;
  assign io_outputMemAddrs_3 = mc_io_axi_outputMemAddrs_3;
  assign io_outputMemAddrValids_0 = mc_io_axi_outputMemAddrValids_0;
  assign io_outputMemAddrValids_1 = mc_io_axi_outputMemAddrValids_1;
  assign io_outputMemAddrValids_2 = mc_io_axi_outputMemAddrValids_2;
  assign io_outputMemAddrValids_3 = mc_io_axi_outputMemAddrValids_3;
  assign io_outputMemAddrLens_0 = mc_io_axi_outputMemAddrLens_0;
  assign io_outputMemAddrLens_1 = mc_io_axi_outputMemAddrLens_1;
  assign io_outputMemAddrLens_2 = mc_io_axi_outputMemAddrLens_2;
  assign io_outputMemAddrLens_3 = mc_io_axi_outputMemAddrLens_3;
  assign io_outputMemAddrIds_0 = mc_io_axi_outputMemAddrIds_0;
  assign io_outputMemAddrIds_1 = mc_io_axi_outputMemAddrIds_1;
  assign io_outputMemAddrIds_2 = mc_io_axi_outputMemAddrIds_2;
  assign io_outputMemAddrIds_3 = mc_io_axi_outputMemAddrIds_3;
  assign io_outputMemBlocks_0 = mc_io_axi_outputMemBlocks_0;
  assign io_outputMemBlocks_1 = mc_io_axi_outputMemBlocks_1;
  assign io_outputMemBlocks_2 = mc_io_axi_outputMemBlocks_2;
  assign io_outputMemBlocks_3 = mc_io_axi_outputMemBlocks_3;
  assign io_outputMemBlockValids_0 = mc_io_axi_outputMemBlockValids_0;
  assign io_outputMemBlockValids_1 = mc_io_axi_outputMemBlockValids_1;
  assign io_outputMemBlockValids_2 = mc_io_axi_outputMemBlockValids_2;
  assign io_outputMemBlockValids_3 = mc_io_axi_outputMemBlockValids_3;
  assign io_outputMemBlockLasts_0 = mc_io_axi_outputMemBlockLasts_0;
  assign io_outputMemBlockLasts_1 = mc_io_axi_outputMemBlockLasts_1;
  assign io_outputMemBlockLasts_2 = mc_io_axi_outputMemBlockLasts_2;
  assign io_outputMemBlockLasts_3 = mc_io_axi_outputMemBlockLasts_3;
  assign io_finished = mc_io_axi_finished;
  assign mc_io_axi_inputMemAddrReadys_0 = io_inputMemAddrReadys_0;
  assign mc_io_axi_inputMemAddrReadys_1 = io_inputMemAddrReadys_1;
  assign mc_io_axi_inputMemAddrReadys_2 = io_inputMemAddrReadys_2;
  assign mc_io_axi_inputMemAddrReadys_3 = io_inputMemAddrReadys_3;
  assign mc_io_axi_inputMemBlocks_0 = io_inputMemBlocks_0;
  assign mc_io_axi_inputMemBlocks_1 = io_inputMemBlocks_1;
  assign mc_io_axi_inputMemBlocks_2 = io_inputMemBlocks_2;
  assign mc_io_axi_inputMemBlocks_3 = io_inputMemBlocks_3;
  assign mc_io_axi_inputMemBlockValids_0 = io_inputMemBlockValids_0;
  assign mc_io_axi_inputMemBlockValids_1 = io_inputMemBlockValids_1;
  assign mc_io_axi_inputMemBlockValids_2 = io_inputMemBlockValids_2;
  assign mc_io_axi_inputMemBlockValids_3 = io_inputMemBlockValids_3;
  assign mc_io_axi_outputMemAddrReadys_0 = io_outputMemAddrReadys_0;
  assign mc_io_axi_outputMemAddrReadys_1 = io_outputMemAddrReadys_1;
  assign mc_io_axi_outputMemAddrReadys_2 = io_outputMemAddrReadys_2;
  assign mc_io_axi_outputMemAddrReadys_3 = io_outputMemAddrReadys_3;
  assign mc_io_axi_outputMemBlockReadys_0 = io_outputMemBlockReadys_0;
  assign mc_io_axi_outputMemBlockReadys_1 = io_outputMemBlockReadys_1;
  assign mc_io_axi_outputMemBlockReadys_2 = io_outputMemBlockReadys_2;
  assign mc_io_axi_outputMemBlockReadys_3 = io_outputMemBlockReadys_3;
  assign mc_io_streamingCores_0_inputMemAddr = StreamingCore_io_inputMemAddr;
  assign mc_io_streamingCores_0_inputMemAddrValid = StreamingCore_io_inputMemAddrValid;
  assign mc_io_streamingCores_0_inputMemAddrsFinished = StreamingCore_io_inputMemAddrsFinished;
  assign mc_io_streamingCores_0_outputMemAddr = StreamingCore_io_outputMemAddr;
  assign mc_io_streamingCores_0_outputMemAddrValid = StreamingCore_io_outputMemAddrValid;
  assign mc_io_streamingCores_0_outputMemBlock = StreamingCore_io_outputMemBlock;
  assign mc_io_streamingCores_0_outputMemIdx = StreamingCore_io_outputMemIdx;
  assign mc_io_streamingCores_0_outputMemBlockValid = StreamingCore_io_outputMemBlockValid;
  assign mc_io_streamingCores_0_outputFinished = StreamingCore_io_outputFinished;
  assign mc_io_streamingCores_1_inputMemAddr = StreamingCore_1_io_inputMemAddr;
  assign mc_io_streamingCores_1_inputMemAddrValid = StreamingCore_1_io_inputMemAddrValid;
  assign mc_io_streamingCores_1_inputMemAddrsFinished = StreamingCore_1_io_inputMemAddrsFinished;
  assign mc_io_streamingCores_1_outputMemAddr = StreamingCore_1_io_outputMemAddr;
  assign mc_io_streamingCores_1_outputMemAddrValid = StreamingCore_1_io_outputMemAddrValid;
  assign mc_io_streamingCores_1_outputMemBlock = StreamingCore_1_io_outputMemBlock;
  assign mc_io_streamingCores_1_outputMemIdx = StreamingCore_1_io_outputMemIdx;
  assign mc_io_streamingCores_1_outputMemBlockValid = StreamingCore_1_io_outputMemBlockValid;
  assign mc_io_streamingCores_1_outputFinished = StreamingCore_1_io_outputFinished;
  assign mc_io_streamingCores_2_inputMemAddr = StreamingCore_2_io_inputMemAddr;
  assign mc_io_streamingCores_2_inputMemAddrValid = StreamingCore_2_io_inputMemAddrValid;
  assign mc_io_streamingCores_2_inputMemAddrsFinished = StreamingCore_2_io_inputMemAddrsFinished;
  assign mc_io_streamingCores_2_outputMemAddr = StreamingCore_2_io_outputMemAddr;
  assign mc_io_streamingCores_2_outputMemAddrValid = StreamingCore_2_io_outputMemAddrValid;
  assign mc_io_streamingCores_2_outputMemBlock = StreamingCore_2_io_outputMemBlock;
  assign mc_io_streamingCores_2_outputMemIdx = StreamingCore_2_io_outputMemIdx;
  assign mc_io_streamingCores_2_outputMemBlockValid = StreamingCore_2_io_outputMemBlockValid;
  assign mc_io_streamingCores_2_outputFinished = StreamingCore_2_io_outputFinished;
  assign mc_io_streamingCores_3_inputMemAddr = StreamingCore_3_io_inputMemAddr;
  assign mc_io_streamingCores_3_inputMemAddrValid = StreamingCore_3_io_inputMemAddrValid;
  assign mc_io_streamingCores_3_inputMemAddrsFinished = StreamingCore_3_io_inputMemAddrsFinished;
  assign mc_io_streamingCores_3_outputMemAddr = StreamingCore_3_io_outputMemAddr;
  assign mc_io_streamingCores_3_outputMemAddrValid = StreamingCore_3_io_outputMemAddrValid;
  assign mc_io_streamingCores_3_outputMemBlock = StreamingCore_3_io_outputMemBlock;
  assign mc_io_streamingCores_3_outputMemIdx = StreamingCore_3_io_outputMemIdx;
  assign mc_io_streamingCores_3_outputMemBlockValid = StreamingCore_3_io_outputMemBlockValid;
  assign mc_io_streamingCores_3_outputFinished = StreamingCore_3_io_outputFinished;
  assign mc_clock = clock;
  assign mc_reset = reset;
  assign StreamingCore_io_metadataPtr = mc_io_streamingCores_0_metadataPtr;
  assign StreamingCore_io_inputMemBlock = mc_io_streamingCores_0_inputMemBlock;
  assign StreamingCore_io_inputMemIdx = mc_io_streamingCores_0_inputMemIdx;
  assign StreamingCore_io_inputMemBlockValid = mc_io_streamingCores_0_inputMemBlockValid;
  assign StreamingCore_io_outputMemAddrReady = mc_io_streamingCores_0_outputMemAddrReady;
  assign StreamingCore_clock = clock;
  assign StreamingCore_reset = reset;
  assign StreamingCore_1_io_metadataPtr = mc_io_streamingCores_1_metadataPtr;
  assign StreamingCore_1_io_inputMemBlock = mc_io_streamingCores_1_inputMemBlock;
  assign StreamingCore_1_io_inputMemIdx = mc_io_streamingCores_1_inputMemIdx;
  assign StreamingCore_1_io_inputMemBlockValid = mc_io_streamingCores_1_inputMemBlockValid;
  assign StreamingCore_1_io_outputMemAddrReady = mc_io_streamingCores_1_outputMemAddrReady;
  assign StreamingCore_1_clock = clock;
  assign StreamingCore_1_reset = reset;
  assign StreamingCore_2_io_metadataPtr = mc_io_streamingCores_2_metadataPtr;
  assign StreamingCore_2_io_inputMemBlock = mc_io_streamingCores_2_inputMemBlock;
  assign StreamingCore_2_io_inputMemIdx = mc_io_streamingCores_2_inputMemIdx;
  assign StreamingCore_2_io_inputMemBlockValid = mc_io_streamingCores_2_inputMemBlockValid;
  assign StreamingCore_2_io_outputMemAddrReady = mc_io_streamingCores_2_outputMemAddrReady;
  assign StreamingCore_2_clock = clock;
  assign StreamingCore_2_reset = reset;
  assign StreamingCore_3_io_metadataPtr = mc_io_streamingCores_3_metadataPtr;
  assign StreamingCore_3_io_inputMemBlock = mc_io_streamingCores_3_inputMemBlock;
  assign StreamingCore_3_io_inputMemIdx = mc_io_streamingCores_3_inputMemIdx;
  assign StreamingCore_3_io_inputMemBlockValid = mc_io_streamingCores_3_inputMemBlockValid;
  assign StreamingCore_3_io_outputMemAddrReady = mc_io_streamingCores_3_outputMemAddrReady;
  assign StreamingCore_3_clock = clock;
  assign StreamingCore_3_reset = reset;
endmodule
